`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OuLqZJQvBwP1fDb5T5S92OX4OOx9UnjIx/usTgfioej1RuGitQKxV+6G44/5K6uXJk5IepxXBJK2
5UXhWk+N5g==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kf/u2ZcH3eks5c2ZTnBo8lBw9GIMM1HSi//QcvSiVCmb+gvpfEarz07pZdv8pnJYrSn6AmsAMoZU
cbCKDDY+9uR0hLy8BhhEFsG0KXNtM51Qn7Rej3gkdSRLc14phs1AeY6p2TwDzdx20hhMRpEc1zHf
1601Agcuv4VGsUZJb44=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gCAMZ8dRLVqKW6HXYzHKBOuuV5+bHoLtKdBZ4aj71oZ08rqyMvwGaTkGDlepRyou4lbos4Sf2R8V
RMl/WaKrbRQqBADwqjYnllwH6pLsPPj53ofpIlPP5bAyPp24HDr/lR2EPUypFudOahzJVUa4gztV
a4Z44ZL5AP/0BYq1cupnhG5lVYt/ozc7RZSabL9XJBtOl3NeXxlHio0+7ikuDKxjvul10su3KhlF
fSWBIznXqLgjJa9vbvop8kvvZUazb653hdy9X1Yg4TUKbY5oRmdMx0CQ07tkf8+gGMc/5UyTqKdi
M/41cefQZFU7ids/DDZ0E3E2vHZHRaSIiyfWfQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cmcyA5DrdFR+Uw+L7nvOCnhRmFccdEdIS2b5dgSFlzFhoSOnIrFAjpUP/XBuqFcV6fPMbF0fp+b9
/aRWSe426CXDWdYbx8uRuCrV1NA8CNYLJqu1GCm5TZT/m9YCRV+/xOCQXQqIlG+mD5h5+s+d6XVC
CzzsOofJO9P07PCN8fIqQWvA7qpwGI7xOsGWNMXo0stNEHcCcNDj5mBN12rdKESpcyICx59Lrmvn
fWO7F1xByl2w7J0+ftpbP/31nmM4l/RnXtytHgZbmyH5O4Y2CZqc4zGlz7zva9n7xCaMvuN1Uagm
FSwVwspzz24/d4yJEv6axJUUyoT+9gs6u+ApwA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fgffjy4IF5gDMhZhArY8sP6iSO/Ck4ZmLQDVFuQteumGgNb39gepsp98PXLNq8IRBGYWHmNvXu+9
ewpjg/E7Qrl9RO0rj0RhN3cgOJz+l3MlusiF9mofV9W72uTr8O6m6vS//YIFferGaDUPrag55C4e
+dWo0Hb/vO3HUPXDDbpvtGe6UpMBjPQ7nwACoJAzI2WV5OEVcYEQki/6t0pSAyIrJzyb7HSR+htn
m8UsZc7TJ/Hu7uX+Dh033kFFuczsxZbUuCxvoM1yK7+C0DLt8FjiaOMzxdc/V7hRs3rA8k7kPX7H
eLSVWtrR0l2q5FHYu5gPItzA0L1OOSMpcuEwhA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VRo7Efb7GH551/T9DNDm5iarjMczbIROhimhX82E9cbFXEDIGfRsdwfoDmDlqltTiJ7Kes8IvntP
xgp/97ae7JHFhCF2QBqJ2e/a3KhdHm3az/zqKBDENd86HsXrZGxQAmxmTvBJp2BVDLHZSNhOy2Kh
opQF6kX0hA84ITy1BZ0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QAg7Bi8l4USBSGMT4MDNYHxF4kfhK5gus1lphOe2yNyQy4BcsprF3Yt2O6H/XQAQCzdpDJtHGFGM
0cCzLybSRfFgsgHO8SeuaDNXg5w67mjkh5HvBTpBTdijfoKiTPCcG76iThkguhQ8EDDlK8y0tmOR
Ptw2b2CQxyGoQSFsCGTef3Ph+1escOPV5nMQRz0xzlKWHJVkWRf9DIuHoMTkQ7y4ht0hNVry2HyM
FUZ83UAye4PORrLGkYoVguP6fxosdDumzPUP1paQoc0G8kSlyHBtvVQHmTNJSFN/0Hkvn/eApBis
hIpAUclDIPcoopOebSTYJpQj20b3X6KEaFgSRg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6400)
`protect data_block
e+UVkPtAam+7HjTBfVAWV8edsrXqg5dfApoa1xR2xmuMUz+8pwHfh+iH/Lo5R5I+MeqnSv7lgtU8
3OOCA5JjQ2FK9JA7qLYJiNkgYkhJuSDQ3kGBoi6vNk0ugPUlPIPDDGnKDe57lqVwUFt7LKaZSOat
lXhdJ8yaJa9eCiMhJw8zPytJcFWAYyX5QUgN8CVSHouXj/rn9c4DsDaZrTEotixHW2QTcSciyRLO
Tm3Z2gVvmtthABfUP572ryqqqyjZvl+jgjiKsZENrkaVk7/ICYR382Z7Efrn+JqKE6kLeanTc3AJ
/F0DNE7hrLLKtxqthqB230hNrdsbyS4NFAJFNVm4qG4+QC0KnmPw3N7HV4+IGARhT7nIGlF0YCg7
oGnrxmD+8D1QWuBZqF6IV8mnobnUN6RW5R2wzsEMxp6lbZGvQBhoEXibCSoLwey7SLlocYiXzBIE
K/sfAal6Rnh+3Wn6UhrgJ8bKIUls+9bCkfrZBm5u5+Pyj7IRHaA2Ot0hlTAjKJ8HG/rWdeFAL4ho
snFD4d5AjxFzh8N4gWe1AUdsXAH9rVaS17RVT9abCpRyLzrVT/fSWBNe2KuzOLk2FO3uYyQHOL7f
BO3wxWwujqTwpplFhK5+TlPe0/lKZih2PXewNU/ElWzlujUFo12anZ49a2qe4HtmbmeqKoclb9/F
o7mR6KuJegyFdAgYv/E+e24fwI8EV+LrXt2icGL57/BryR//4XFTxkVzuD7p9Q3c7FwCt9+HIh4R
PdAY7FlkK01oKc0V5R/ENknXLDaHKIUdO+vbqTzaX+ORGm4PBlk5FzPvcN/9ULH0NlqQqt+TD69L
JL24KynxzfYTHyukS4/B+71R5DH6AghHj7PRpRugjywz5W70l9q7SNyl+FPZLGc8OqDEkm0Uauxq
DMzn0wwr+uLKplZuH9kRfaEPKRMaoGyD+hHyBpf7tUMIHPS+/d53zEtRxRZ7Y1NNZxVkZZjR0sxd
Cp2Vhm+w62y14oa+4/bE4NWIPkqL3ZUX2dRuHonS9eKXaBdCDYEVRg0eyJVcXEhYess5gcFiAB0q
/7Mt/eLlKinPfno+x0One8U7178QtAeemJYDkrjBwt3ySHOTKGGYuom1yCQC/p/FclCqJgH+XNP5
bJZWc3ekwvYM2D+X0mWR01ezwdySSr+p0Y5j444OO4Owef3/yN+B5WTzy9E47pqYfpLbJAcFgVQE
Epi7919T9iIIAlskLWk1WiDVJ7cuWiT5OUalZ70J78P/ORH/N5tVAut5AGK1FhXkOr0ctLDaKfU1
IByeCQGtOBce6WT/FOhtLJOe8aAtYYeNPkljNZ8Vsbom86jMCt7Atsr2rqxucSxgXxJmJsBKAUMf
/82KJoZJoM1eFDfnzg6GF9mJvG1dss2FznlnhzsCXdeEMOiwshzN6iV8o7kRtAFm4TQvS6104vtA
ATsfwQ57KWDPoPE3K8KQAQPU8ZeNhdO5KrLnUGHjoegWo2O7PCgbnHwXnx9pWmi0QQ/cvc1edoxO
1pqAtu1L5+K/rMUc7mNKU803pMiED6b1tpiKAfgrF0r9u0BZHcLjUbhHJIJXF4LQYTETjrB6iJEM
F1NvyfNGPy/Qb4tz44wPBA3C69Vd/zWAOpKO/CMV7U2Y5YjM1T/nhF2vnklHYETtj4xJxDUX73Ir
GmGVFYgEnex3h496z3I/MM8MYhwPbmap79UOXp0pwcR7T4kp44zfUaPU5uZqkl/+xu598IiOB16h
+FO0iz6KfHA/Ni2JQcfqJ+iqMT2VX2dfeQzYmQbVxuKAENyRNNSZX//GbJmI3rpbzaDkEB8UrTho
Hzp33K1JlwSMMp/xjCWHuO5XW1xm7gXnSK9i3gbVUY69TV7erFdbpZukkqnCcz7jYvx2x3QReYed
QR1lZnrY6tp34K1Z4xWWkEgXgHoVRZeBz4nwwGmDJgMwWx1a5l8RPDq8Wu7zAs0+kPrfAlm5ySKQ
V+Ry3jH9CjDFgPbfFdTKAR5mZnYI86JBdrY/RjfDzr2F750pp7Ls9bihmui/qwqvFKH/6x9jsgn0
xpoV18BIHgNjVT3adpNDMLoRMLpiYWiaN8HZ1Xsvwr3fAPR+GW8+ojwexmHYSNI3i+v3n9JOcFpa
9OvHdliryuvI8Y9GQq/BgcrrhLDR7GbPPLSYpDqrUQJF6Lb4LIjTYAPPDiN0q/euFfmK5MpEC2vD
TRNaqG5NrVC/B0noedLq3ett58YXqcv+8oW9HX4NeflaDfUtzGvgiYr0AiUPX/xBiUaUrgonO+qZ
jWxyUa+NiolYby0J5G7bu8WkNzGe2it524crVVq39DYKInv4X8nn4fFi4+3TU+jKx4s0RGUjfc4/
yeg1+KJDmDVSIhzZp0jxaFTDK+NJRLOJQcVak6XAlWqiaKKeeN6Nqdo/P6szxtykqfJeX5DTUG3z
f0GdStzz5OUL4VpPw7gcGNcbGzXcJMwq29RLo8tfUR9k4A5zuXhYrVCDk4dx0BeqA+3I/pE8v4qi
042XiW6DnGtJ7Mu43abfnBEAgyguy3GZ9k9fUr1NR2OZT6bQU4nrTLrWas/CF5q130STMTQAihQQ
36qzBeUS2bGeqsSxKPZxwO03kKI8h6TESAk8i3SCuNilKjzmZtR99o7xPosQi5FpoPcVtfTiqoTw
+Ty2kbLVqGtf18Ozz5RMWXFpch1PXVdIFeIdhbNwsextuJlELIoi0/q0DVHO+8uWjMsTKwudHsxp
p73VncP7g0yN5yuryylBZ4Q4ERs7LceWBqi9DnOkW58JqbfWyOq6Z3KVHzTYlkrrLC3jo3q3IfVF
y1UzLgJf+2T/PJ7qNhJnGCS88yIdP0Z//3Ip8Gl2Yl1jB4H8edtxyyGf+XQYad5SraJ65YqcJXny
Wc0dec0UjbEIfM8uivMyxmWscg8gSq8NAC8vnvbjcqMqaoT0Q4sa/JVbHYbXCkO2G7wKroGAS+HW
JfBfQibuasn+TrpAvw2Tl9DqWZNw5DRt9weDKfAQ/wqKA3vjRjfsHD4dohpzkpgLYEVpoOy8IqaS
JW66xQlWeKGGVe7Wu/PzKuzX0l7iiQjL7nVavxAKSQPSXor6UoxuBsDjRfA3qxYE+QdXKkHo0+h6
6BxqkqELQ32i4abbHK5dmnkk0m8NeT/69G1WCSaeBN3E31qJAYdyF/Y58gIVni6tkqSkc0lJwLL6
7rxXtoF+oWROf4QBro6aBf8jSTHdkbF/khnwxUSOv5cgcgNY58DaBmVgCYYHcVOcg4BmVFx/hYDG
/zyhWjDn4OSwkFE5hHYPVwbNbYZfInxFAurY1plU56oLoq+fvOltpDnHhPLQjGfRNX3ij5AHVn25
1isqlTte4yEwBvE7SxMYGHk8Qh9PQoEAJC9vDfrQ3bajrSEAagUgfph5R3lL6ryBB/UqxRnEGvxA
lT1hBW3qXvSN/UGbGACkBNkA5MccKrvzY9x57j9rljcY/V1LR/ENyU6zzwnHDM1zo13CrbWH7h+t
APNVJ7YCjaO40z43ZPVvagPpC6wI1o8SImzrw8c854H4I4Dv3LzhyjlXToxHXOoYtS96VFhn4Dig
kawXEJP0pS4HtBPv7iU6TG5ruyD8UZA72wE9a9O9iJdwwgPvNYor5G2ieR9cbjdqZuyQ46EnPq10
9fkSJewBSBqMGV7pT/jIUgn3r5UuOxw3/YbcfhKVFgoQmXgpUUPzHbp94Z9GwS6ad8hpDWred56y
k5VjY26QNoeiJpX5YYNbC67OsbVzk68yPLX5Qwss8A312hg+fV2opqpu6GD26JsuIAQU1f7GUZlx
FfcqN0EM/iWJ944vfd/LG2KJOHqsad9xPbboxJ6RmLty2mJpymQHGZt48MIyexlrAazdmuxmkUz+
Ieut6+fU/7StfmtKeQ5zDLZsQuJMYDZMaWDstNbpk+ZnQoHXMIe5/7ABWi+aUFheBvA/t9jsDF0/
RGjt5mH5g8JCqcb8JJeImeUi2wEc2Ec1gls8C4Ooj36YYswTLIEinw7rj3Xv9HVm45zAOJMa3B4W
Zs9PszCSVP/ZHrzo5n7GeA+BIImPfuJHCpR4d1+i/rf2u42voQnTKkMZKWpvpOFsKlSPlGtmpzu8
MpyuPN/igJL34PqlHwjFC39TG8091P9tbKwa4ZCy/AP+X+vOP/zmvkIk/gf5uBKyLDxw7jEAzsWM
EUk42GsPVKI2QMi9TMI/KxV1sXxgyYPLTVYworlDzgesvLuVvNgjWX/QBaZKRuqrJ5JQWXcPzJLE
sRUNaLJkKJOzXbMMHxEoGO7JPltPzmtixA1rojggjh+lPy+TkRfnMyYbUjEbawAsBDGUQAO6LzD/
x32Am+O0fjdLo+N2HTJBPMbG+rxhqxJunegJggKLV7qF0egcP8dWc90Fm8h6+ErdzSPf4Kzzo/c7
3fVTHXDi+7mLMsmoGxhKKs2DwYrcHj0AFAs4kvVaqi6bwqEg08roHyzDxmS2luXK1GcKlCiAJxbk
W2Nc2qXpimOsDscJ6eC4ymL4gmyp+cxnabtOnSoKVEmGr5aYIWMd7QjFmiRUwtnMZNQoo0/D3zoe
y0Vzkxq9Ol05qLaqMpXGAyfJgxPrje8y1A9YPfzoYBpMrNraQiWMNutYNsRF0IfChjEgtALL/CNh
oXJr7j1LgDotzb4snhyoNOVrSWfs7BYcKounDdzbglOFbhQPbX33kkhqXzN0aWM7rQ9DAc4ebSXn
ipGTvr1ADt89QN1gX9efQJx6bonHvyE4FOBcjidtFX52XHaDtLYZSR3LekLShau5rZHHiMwduvIK
YrzWL488hAt6wBMC6X9hWhuaHnT15oCNTVO2IaLsYDXA50Ognv2oCOWZenWEkTBLI80yDwWxNpiQ
5d54fLEd5ZdLdNm57fG1ttP5Kiq3WUnRGdBEmUIH6SRPRILyDMRnI+S7VIxIsBk6zdvGaOT9N/ad
51HqQudiJYU54ONcdAOQdWrmaC93LHOjrHCO7KxCNGphkVXiCNw+pLic4+DNIV1YNMG5BaK0iQfl
Cl9edB0FSKUO4u0IWbG5bZcRw57jnIUaLqx3yiTcLlHNE2gx7KV4N56P+fCdGfKtIWOW8MHp0fmh
OXlzQVOXJJbysatsk5p2E22Psug0AxhK1CbDBdENor0wEcIex1yiNDczA3Sd6zF96n2Dc1jVrioY
wuW1cKD77Qr5uTLb6r7msXMkTCJIwqAQT+7X4v2hWCyYb6hDrm2gKPjXqUyFEHXs9VORI6skNc7e
/QsPe/aFY8FQcCQmnwt5U//f5yeVHO+FajF56cuXfj3jvno6wS4KxOABsjypNQ85on+0T28PsA8y
MrGYNiawqlWXJHK+7idw0Ic4qxpeVBO6rq/FycSdwi5FCVLq6Q/ULfilmF1ScDkJ1eb3UeE+pDgB
5l7m0jRD1wVjxvjo7cEwJpDpWO+8JB6MY54LMbi0uTP8ijNy9c8Qad6fDU11GVVkIPa/Art/Vxju
AqCXn731hrdlpX8sm78ssb7d6DMA2q+4SfeWSA0tnfgvgCSg/7JkdkabbPImY9ex45EoHQGmdUiC
FVgl58euFr5yw9qe9zmJgRfXWljnPVXcPKjWE4cg2BWwZcGroh5JMWn5ECEEXX0tEWqRhOoWliQ2
BpqFFglBXrpAEd7xRKi1sFfXlPxdmcgrlAs/FTKBtCjgOnVGmJqfw8mHtQmBZyPejbBRvqJI7Xit
kNsmNyYz80X/AAMXrp79gjRyzrZcn5YcgT2Y53jzGW69j9kWTEOkrRUf9OWOT4iWJcfKHgL/wPPh
oCpqLRz1NoGWmmtIarxox5bfAJustDHC1z385aS/GBy+/EinGLRXvYSYW+F0k17vjF/7LTyv5Do8
z9BCU/8kRJeDAyZ/d0HngltefLLfiy2nSrhSLXgMuJtVgR9yn2pkklaSwJbT9S+Zo4zT+AWFcLXd
dJNd5MZ+0t1qIDAjs/fKKEvzRXYlaPFWkJ8x2VNm1kX8h5Qynp02Bpu3MGR3qeovhfZdiQ+/otb5
kVUK9zHjcm6jyBVrD3dlx822sIDCbDLCRoXxi1Z7ocYRJhZXQjVnhLqidiVekaEnBAPzvjxuy8jf
hfJMgz59mgFRe/6oWjsEN3B9iDMxxkA66S8C4Z+4t3KZBShiTyxQ4Jjp1JJEXh4zD53CiiwW3eoW
J0zxN5+EUx+9oSHFZOxm12Ee9lK7KiFNJ0nxEn3sPPrG6Q1GbmhFbNIBespNhrl3dUCodK4IvxvG
tZv6Z57CZgicdSBdcEdX09h1rQYfXY3IvJtNNegXOaxhQiFjLB7OovHNrPjS7njpImGaUjp+m0Cz
dX2onBk4DFVaTABG75utx5YDQyNX4jpi10i+6r1ybgWQUnrHcG1Q3CnB2EpH0wWhBg65bclAUJR0
HSXv7BMRNJCuK6XQfdtFUf9DhOLEwRQSwZ9n6Ix9VGv4y1u1v63AWnqN3VCFPWTVX50A7d3/Pu6i
EBC3gSoIXrehndTaIROPvDwVO5/QFfIS/0zeWaa1ipwfCfbkWqzKp9DiOEo3zLCA3sjrQXWGeX0g
2YK1X8utmZBvpIN1ucy3TXrqW9fKmke1YuhKZtyIN+rQeVC/eYWbUto435/gss87DrU9trz4tNTT
c9Acp/JySQPZn3M4sSoVt9jkv9MMhsMaFOo+KgnBChfhk+nExEgzv2kBPDraoCiDOQdVR2zjE/YR
tgusdTaK756DHTusMVSVyBzrb0m+LyG+ln2TiXwAjbHIsg5vcGnKdmAdSDJ3svYa+u7aQ82n1bJ3
fECq9w9yhVxIJFpWlZWZ16Y5v0P3DEvbcKeT1hI3ylYWtbppievvn5n6pS9kU1bh6hYlgwEn+yDj
OIK8GVNjlzfxlsp4mvhhjzdX8nfNxaAXlrSJk9Nwm0vLKOvTMu4OUXzD3GYnLj9YGfaYjiVqQxKs
fFyAgOzOzVvtDaB+oQ6PiOaKqhiuxyg3qkGpLmyNYVIyNStW2vDi+O76UgrVmA2k4/p2gc37W2s+
bQ6M8NrqMBhujvng5YVDUXAu/Jx6Bqu/wZ1iBscEdQXJ6N7V8i+EOnLq2lcFYkINcAUDcZVEGvyc
zxvreqdDAaa4w+q/5zlk0tEzHCvQY4+VJKnTl5ckrLmnLlxunkTmmzm5CyBvAo2tR9R9q5HL9uij
OiugJbScP0RYii6UIJfblZGvtY0/gxNPhqjur6a2XVBXvJHi7I/dsF1db51YmJtf9gp/JDuAy9Eq
CmyeETr39tKPH+AgScgZJuPGyLM0RsYvvrj3STX3hUBNakz8IkXVQqGGxL5AVwn/fCxFCay1nl11
L59oNR/rIftWe4bwhzJd2iUqGL8+t3LwB4USubBj5VQDp7qyTKkWduuHhjUV3iCiudXZCzPQCifb
mm6gDWXRgjnYmiG0urtEzyx9KmtewDnEfoguP7mLZxeMn5bAM0QwHN+yukIITuk5tt3xLoQiPTdD
itn71hmr0AeLPpeDivzVw99Hko2t/se7Vu+DvFJR7tAf45X7eNLtVVhF586RlOmOwRoKnbz1pnzi
r97wY4DISQ7G85mUCzsia3vmCcnWG7MjT+SKKKprg1sIn7MojRY/yJo1TQyaxOE9V81Zu2KdSuXi
0SeRV9cNXn6l1aX/NOaLttxPOmsQ9YOdggmJOl1I70YCqhe4lXWk5RGzCZ5XsXor3AX9ztQYv7Ve
B3iy+uw75D4VZsobRagErv2apbfRwJVfOA0RdoJD8yOi+aJQIhEIzQoY7brGoMWGLHHmKBfV3I41
LoZJIazS00t0s8FwxLmKh2/Xi2faSkQMHrHDmPQu6GDhlN3X3qJTXcBIM5Py8qzweoOaWOmmcKhy
3gyVJRjQs5kJCKRCFt1YNE52qwIk/zUEME80BmMksoypE5V2pxnbxAog17Zc+a4AerXhZiEy+iof
hGZxKa+slwyXrBLVsh40hnTmj6+lsMTOfBLZL2jZQBeUI9Uv/hOcyXKtsSIWP4JhIRaXniPSOvEQ
nXgWtAjQX5DmDeMQSG6fLoLiV3vflQwCZBYf2/gHschnl9/X1V4EFn6CwezUNNyj4QRhwI6J3+Rx
wLeHimfAuMzTCea/Hf61WIQPnxfrcDnPIGQmtpm8GFztxdZ5mMfleIb66LT4by7caLpeKuPkC9LV
soo3tfmXdOEcZkMFMxHfsGx9JPSPsz3oIOccqFx9kFwb6Xbiq5PRom5y7pquv1k477qIEzhqT1mT
pBogLX6S+2gUo8eECbEGVE7ezEuOUkFxemXc6cp4v3GtK/2ki3yXWB0aRloaKZgVJldBivYRqV/K
xS6MgOPr2ss/bU2wOr4s+WU2TsyOWS+p0QvDJ/BP5nYdpveHXO9XSrrU61vI6MXlUmCuIZ8M0NHd
kB1Uiq9Dw9fJyjUsJYD5Z3Bm3BwWqsazBtd5qa/oKcsPE6yvB/oeTqNayvqQTHnXZt2uB6+h2OhU
4KPEPSEhfXFp8QnnXUa6p9OBQ6dSm9k7QtVMC73aylmrpv9QPk0/Mqw63/J9lLCsOMHQn5sTSxiv
tl6sDvYwB1kg4vVL+nmeRA==
`protect end_protected
