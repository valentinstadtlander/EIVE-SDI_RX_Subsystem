`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ENCQi4QKL8B827a+130AYaVwDLF9GgK4vgIJHFnbkoR6XRs238yzytR+FlL1pn0FQtaJbcqK15HD
AlEnMa2/+Q==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wGBnCMSDC9UYWmogpnyQZ4rhZ14L9+8yM3O1fn8HVfnJA7E6C7YZ80mH1IZWlHrOibLsDSUgYv/y
0vyQaCDOH1vKm5cOfNcdZFvipMt895dwisvWqB9/Fq//Vd+LWoGk6WNa8h09b6UWY8kNEU3qzkDf
todQySflBE88Q67E9xw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OtB4hzBWJNqRnuvMXfJPbrLcLA6o35Iwahh+FCEmuT76QPHlwcN6J4mZZ0R2KwLw6+aOYsWzgBZ4
B26gfW9L6W3d+u5O4oc6vKtPulbm487YUEU3TsjoVRLukF8IzCK6tLWIN9untuIzkQuY2+p2F9Y7
yCNli6o+BbFOwHrPGe9aXJc0qr2iNAwEgkv2E/xAwpZ5ZCN60t+NsHjM9K67CHYHbYFY7m1W1qlx
47+WNnQPY7DugZVvKPHIGA61BXl7xU8WKwWwxr+/OF1RcVwqYfUKApFVbzFknhl6hQR8+4G+MBXW
w+m+D5oFwroI+L19LrmeYfBoYTRLcpc3DUsfVA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O8ZCkpN9JhiyIY1a0d3AJx54naBKOptXKrE4lcqwyox2ndKm8PLvOJcg4nWV9NXKlekfDdk4tL81
V20waXH0jE+NYkHrktqxYdqhOlJ61P2eai1GtUjzBuNB+DPO4qIZecZPll2nGyZcGSL2vRjyGJaa
fg82CQ3AmUSk0PsLVNk7io2lMy4AqqvfDt/0SzEUzitzgwGuA9XXDiPLE0gbF60nbwGXCALqnodZ
tirNeZbQC+klhHYBQ3Ifdh3QswZ4Hi/WqqL8aVZDJ90Rady6ywBGgIiURX3ov0fPW54k8GtOGbA7
J4A3TxhUduwZNCblq2uwNJHXPQCUc1PPXkeZOQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Xhai3q3GDCAhWlYoIS72fSSzC+Yyszz8RSYZ7dYEK8qbx4CpLG1MgwS2bRFYctHSMStV8dqk6vUd
ItFIFLhlpmeG6EJOQhY0WPOMR9+fc9xJwAwhJkwPQ9j3/fmr1wmvJI1IfaewNctH+Adjmd5X37nZ
vC1pf14QEU2i4cIsR88SEfaJoysWjv3eQWvadP5qT6pew+sl+1uUtcvOptB1/qZrzmj34A2jTQpO
bhh7O0RarZ18QWxN3SZuStK9IfDBYBfzG/qDQpyiBjOe1rg9grieRRFHzSt3DukDkH9TTMlCeOmm
fNvsIh7340EECR8zch/So4OMqEG79L2woXe3VQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uLSLTu3VBhGpA1V/h+KH62bZ0BVT7b8vYTsVSj3BgonE1lZjzDPowPkKuZg2EzU6H29AczNI8cyN
t++Bohe5w5EVLgMEJaAc40xuIFDk3Tldf5Uk14g2X9Z6j3GdHltlcST0jPhJUsn2WTlKN51Mnn9e
XMUEo6GBPLdTmkKIu6s=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UNpYg+L7Qzt0LKrx3l2iiraYW2BHKDRXamwKI/ieuIcQ2/Zvyd55tDoqGMjGdpu8S5lG0Xl8dgv7
SsHFQL3Q89vCC0eqTfYFZyLyGfnqi18CO3R3Zti7nX5y7cSxKAzYWPf2n/3Dhr59jjFBpde/gs8T
29zGnAml2VdJspQVkqIh7J/UaZUPKwfPggSd8cwOU4LPNJEUQmUTwYoya6sElpwdbu+wjb26AY36
zai2UPAux9NcmWDXUp0vF4fchM4eSpv5h8aFNCbwjaKUtB28B67f+6aug/3DWMn4opUwLQRrcMbh
ZYNFyPz/lOXbDmWQ2mhQ1lahMW634eujd+vjiA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 85808)
`protect data_block
HGOR8XyKmx6sX7+05r7EaO9WSTtfWubpEvdivXLnsE9g3gjBxFEp1WrBGmZ5u10ChE1i/J68gQh3
ZgGZlXb92ix07qUsu3AMcL7IeQdILydJMCb1Rq45e2dT7MDZ28Qe+aCqtpMlQvEWOd7p/4nMyhp0
n4H2bUWwD/BQP0jfeEo+1j3vWM00F+2FqbzVm38ZoZTSBdCyLEGYLgxbzb7FYutxqPb+3G9fnLQO
k4mrPGL2TPm0U7nNcTf3GZhm892il18z/ckFBI1LHVsfRL+C+1Up30rTQ1Ja4luhDD0MsczHLPCP
9e6WJ1s41nPpfOqrqxgITYfd5IW3EU29hq1NQWDXKYntjlIX0jlA/HqTOR5eL0MMz5DWnptTprUZ
T567UkOOOnu3vPdQZPcwaPNsCurlhKUkJkYFFvJXlDRGwPhjdZ9ESXeOzPggxGT6TaejPOYOqm/b
skHLr4yz1lkC0w/Ehj6R5sf5LMl5UiINdQNsEaIr3CFpdqgz0lx9Hg2LVKvF2Ta3PV1GX0stz+Pv
SiU9XauyYchLSVQjqKzLhKPxozXy6VKkSKcbeVRyq8/n89SoK7e1VpK7HBWICfNUBA2KHGKDu8Wh
m6JNa2bruLLJ097fs1ItZN+RcZy+dJspzKRHxlzmfVrNxt4YWH/iig1FHf+sp9bvsm0wbtcP2Dt/
1oixSQakbP5t5vk1qfDvv6Vw1M+vVUGFtkyr2e+tTnJhx+ttN0hTxDjCspOZXFQlRnULbw4K/MXZ
/CwoPZIKH4KatY0AtZdy0S7+GoDuzMdLciFd0wvYf04D3pSzPhpmvVWEV5lkbbHVjD9g4hXFJ0id
Q9A45LwwfFx6hup0Zy5fGZuliVAYxKvG+ibIoELosLFaCzflAxQDjmbx2CCYWG7BFotLdmqTTjAM
dCa0Ey4cJ8QEJbFOyMKgjqFExwZx/Ny8/ii+1jZvl2lbQSy0I00EVtRRy8Gemky0jTTHi7xN5Jz5
7K+s2rRVJD+HuyMkdIf3fl909kkBo86QHZZw7xe8QI5wKCdRmNY0kY/dVJ6ZSLBzNVNjnlVna4I+
Q3dqcd/1JK9Uc0MHPQI/lXJxJ7XwXS6cN/NQULXuQW5/WQED3hCY5U6NXMdguw2hNps3wmvdQIjZ
8fFbiHkKgE3y1HnMhV4KhH7OiYpCbqT3RlInad/Oh9tB/gQitUPTipQX4q24FCip07g7PKSFvPNQ
MaNlgfyZCl5hQF5Ecw76o3otPp06zeY3FDKX8gYOaUsRz4NSuG1eMv5VvyOQ+fiBYEUy6wLwEUVM
gISsE0lozfjTtj4+wjkTgUWX5IExBkLP22nxYoADuKClYEdNH7a9f58EZNWOpHnuJQCv3/1zdBWf
HlHDlVbHkLEeF57xOrdeU87Dv8Gs1pHhEkrVHLrUrptu9vgKx3LpE2ElWhf0X6RaLjksfXU6lubt
I6E+aR2d8Uc7fi7zxjEyKsCRa5WtQEOoo5H6nD3eYWlPISqHY4dMkE6JdcA1Yrkb9yn/L63A3BBP
xEnkSp/VnRezV59o/uXkE1M+bK5zDMMOnIhgt5C5zIn6w0Rg3JtW+klo7fRikuc4E/CkQ7gdRvyZ
e/50SZgFQZu5zZQe++jwCbpl+qezxil0vbOwouSOEyAymXnpYSOvHGXmX+jeCJkEgKT1Brn8id9M
6KH0kCzSK3RAaOJYcQGtUNoIcVDMkUBuD9L+CIy4+sBPZ/BmDHwJecDUXmjowu5OTtwm9LdqjSyO
whRA1A+hbgte+o1scRHmGcMEqGPYeqB6rCiBZstfZaGDtF46qVOCNaZY1+3lktK87QODxuqlNsJx
yXwG73FLB1nCgKpVCAlEc3Ob8j8lh1ASbKh1om9LvEdnyZUcD65TeuflcWtViq5K42IXAyrqNYAK
0fSEore31/U8/uVD+hfbn8SyQv0LIoo4ApiVliU5q2hDhfDHx6mbinrqQZIRqYPEGfSjqm0c6XEM
OsPxzLBv7b+OK0KNMjmoZRwXUKflr5FUrjgZP01J7MqBZrqXLdx9pNQDxfXsem693RNYkpGRWha3
o1CYXU4fQ8V7SlT5hXFgMK2LJCAVgpz6NKAFcrSiqxRbgZguhT/5WthtI/lLO91QEAh56Ho5J7NT
IBtDGgwenkCz7ZJva8Gnl8Puzvq++3OTHi7Z7U9TJ0SXoVe3QCA23rLjw6yLcFLY0/phN+h0Dc8K
InWY2wjxgwp/mCh0Mhf8kv0+KtOAlwXkRVenbCN/vlmzwOIVeAsIIgI+6PPvdX8A6FchRgzh4OTZ
WwYV9EnAao8jV8pa8NY7gz6xjup/dx1YFlpoKvkkmqUz5aTfzQJjfh8ljFu4VAeLP9jFcAanxMKs
a8BMnhD6hKzHRovAIN4M2owXJaJMq+kwtQfLFx6i7tKWti+0ZJZr6dWg50rEw+3bW0QZvvTPcI4I
BRBoJnCRPwnT37VxZUWSGlfA00ugUR0nZPdJY+d7sAhlgY3dsW2rTb/6V/uE8bnw4U2vLC7zbpdM
Nf/gRskHLgX5L9O/8FMwdUOewoCveqQAZpu+sTHWLvq2oGxERvj1W8kII5gyjx+FK3du84mpKkUp
i1WyclY+LjkWyh/lX2KOMkBHCPuvyBRLpqS0Iw8h1fCl+JB/I7EQs7E7VZpNNYXs0tXgztmkmo+H
M6Lu1J9p5YX8f9m6Hyc70UOqVIDazImQc1xi3FfS3KJu70uvDG8P9nBrHNvse+ShPTAtUVYUHweP
QzgL6z5gQk7cd1J1l2gBNC2+Ph35hCjX4ykfYhMWVnRzq0wAIFrEcAeEuF82L3RyDxOPcU1StaKD
zDS0OLw2Mg5G50g7sp513MraJItHRFJdfCl2O/c2Y0NOL8UYXcXa6AM72DJeFHA/XMVYROcmYRJE
SlBiCqJ87UF9VJlfSM7/rcJyM65F5VkUK+QqNRS6mjKkzcNmmm7OLOckVmatrIlSOtN8DCwqg7zV
HiWy085CvqpcAcSq8mCt6EWoM/S6PmUnx/1G8t5AtDUg5f8wperDKoKiR5ldGHie4yQuW0640SbQ
oC8iYfvIIEtkpGqFZuAtztxY0dhGu+VxkuqXEvFXdKGsUDwAgV3tUeOjo4ZMsCoSrLjsBVgXRgGe
1KE7/cAG4Gc6PH748srU8GVp4S5z+C6ppVdaxdJjpLMIhP0HW6/DkLDrkljBeJUjp3pkwg8QUqb7
bs/tjelMA3e7WPTSpDpweawV6f/zNzaP4Q+HP8NZ038MbuEAWhcFQ7E5lodsHblAV/FaZaFLA5CC
6NwC/4t3GPsI+V92VnaFcVoLb879cAKy57+h/gz8TT09MnY1YOIYHg3PWbeCHzVfka17QM3RnfXE
neX1PVmZQSpzUPmmvOCEBO0EmQSm+j9fa7xK5Ho9Ohr8TGgF14O/1GQtzIji4m+pSK5NSf5owp3i
JHki7PT52e//EXNOdQVQDwlrPLYr0B62TRdGJ/BdCfidxeoRJljYr59fQroIHnqCR09+Q9U1ylMr
KSqvaDkdjSAw/r/swOLnnK0bPFndH1NBSTQvmM/U+aFK9ESal7z9qldKWB2+t0lJQrZ+pPkAH+nE
lZz8rDI4HDD1BxAvMK4i3LzAY5y0ew80jctz+vj7AOundUax77ptMgq5wJFnRc+U4lRGuqJylh6Q
67B5ZS0Cxelli1rUNUFjqIJa1rN41BShAF1w0L6PGusr+W8gfBW+JCE1ZfGoG6UkV63iHvrUpr8d
Qnl+g6rUdss4BuikgQeO9eV8RFEjZNkWu6JpkW/PcRegSdlTUypQlG+oroPAuDtYAyKVuqiL1hUL
kchrJjQ5kJHqN4gwnLN0BpPiQztnOKM4zgmPZj54eGCX4MYkTA0/G+gdDhFyAX+c6BRvJ0l2QMRh
BhOeMy0mDYGMrfQWNRCuEXb/nFsRlE0H/99/PyalpayyHqcYYWTXW9lbXE96vwCclcdW7M+pgoxO
EzftW8rXMNhG58Kv6cDpKnCBoUtJsjaVTPmdsdCzFY/M9I4wIU/HU8LRsuiSShRMlvjz1uPE1BZR
VjrenATuEzqmC+NS5SJ2ln2tjKQCZsEDt8tBlQfH62SmosrZ+zu50T+CkJBnMWJB7ark40vYM0e8
0pwkKuSWu3A67ks8RhXjUJw3lHE7ngyN8A7qI0gXvf5E+dThOAPT9uaK/LJvyZtWVB9XTK+9c/ck
5mc2q3vdZFbGy4XIBVvn0jcGT4KSJlHpDbTECNZh2r+mU4pqXMOUkdBFpnzGk3ZidnVOZoyzJi2j
nmRaIbmRke8sN7alKXL5tvuENcBzTgp1oYRNFc1YBzILZzowcx6dArgX9AMIn1vcYUDpYHcaiZuS
Eceprgs4BEqLSwvaXGYEMm1euySJ9XJa+r82eQosMernYy9otvXIuoPULn2pGy82XRk/xhwBltqa
Wn6dabVbbTw2IDq1jBBLDz7QbZik8tnPJEjOuD5Ebeei9eLnB91iSmt9IUGVxN5KuTjEJLZvYA8/
Pu3jnNCXFLEQ/klwIpxdSYA0+Al6FdO2UtRo06Fyh5ZA04WHyAhA3y8idwMV1kgIKaN6SLNEbLHH
pYR/aewVK5X+K2stPOETt59QPhjXljLUUaohApMCDn8nWbn1NYuCEV6zGHlBqTxM4ik8Wa+rHejC
yYljTADc3AQ+9vLmGVm/1FL+rTwa/Nji+aoee/7RqDJvE5CCFKnTovwHG89S2mDBVaKM6e2cau2v
C8yOFbwcGxlvo1BXKIlS6e4GtTrdwP2OqjsxzRbm1TwRdTTs6mUjgmCPczJD+hRzx6zsDf+fT4XQ
7cyH72fYrYB1KSGGKc5H6jYRnaELvMqW4HLbI822tos8pOuN4atXxmfOM7NtexkQwBAMSMJv7lqv
SIwJrz4AkAMRXa1WlbijjA9Xo5BX5f1ean2M51Ys5pWlkRurm61alBglAwc+JMhQ11N50rKl/jtq
akq/38wFL/z5j7U9PeIVBge66fi/oik6oWBDDsroLki8EoSoGlSiYmK3D9V3JVcVuxmPUnI6+oQH
OIi4wCvg9EzcydPWYgqeVTghzmw48FPDMgYKq97eUP6V8ybXtSKAHoTUfFgNSsuAvFj9GkIvdnbk
OJeX69bC5+iRtOVYwjI7clg8uUqX8pFWGhYhSaFYEoxQWY9PsPk2KFrrhA2jLCBquvX2QQZWUQfS
a0NzmY4an8GcHc12Ksb6W4AV1nKJZQ6PDY747k4xelWcFJN0JiPFPWo1KkAUU+02We43Mr8kuEWr
7/QWfAAX9w+7zuTb7X51jVP5C1hKKoE2fKoGnVry22VT3uNUA1DLHdqOTNtGlTdVF2EqtEdzcNz1
JYaAWFkZ7jXN7DHTLUmbZAxmUV1Unx9xPifRVhIqAMJ5agYHLsvFC23mivc70J2uOTEx/ix2bToy
z1YAEOuC+cefwTF5kftmkHSZlF2sfKY6FGWFkrjEGoGdt/nGh39rgnbekgRSRzYOTxUgst7ye1BP
4AI5fV/oQEgDTLGrX9WPu1HIn+GOe5ebQDWsP8SNAIwYH0mo17R/b+I6QsvFxzmVNa0GhfhiG1Ej
JNt3DsOEO25NpV1AHb44Jq8pbiwhZYwkXPqHo3XwQJRzaK9evuwX5Tu8AndA+MHzbTtux2dkAgea
mHkR+4mQklErp8BX8MhWQxl0hDIQmGaPTMkZyz6Cij5vQ37R+G17l/zw9OdggPxL2KlqSVP5I9J+
xICpnDWqEu7p2759JQiwxHRx7zq64kBvJ0qW4NQkz5l68g7eMjYF8ikGLYli/kazisTy1Yq3FXZp
T2P88f7TYmk7LzCbx2b+w8UAYWih3DPcTyY1wEEloAHZH5474qAuUEloCRCT8opBm7mG2Bs9XBGR
lSF8ElaRrIRdj8Sv+Dh5qotaIKyqLaWpil9iQ0qVJmtpHV1+daENOs+ZDQmeYfQyo/YUw5fCj+cE
zFMbgNdRD6L38Gvow1VPVqIFZYzvwz9dnp/QHGQyvcG7WZFyT2bm1eqEVnXI3Rm+FBUTnX6/0wNR
dxHeIdJdH4KIK+0B3EOTx4TmdvZpjfH1l7/HerVovAskBQwzzdTPrpVXC0EjA0m5taASmyY6u5Sn
gcVnmVXKwSsc5YPbC4UOrBYPNrh1y9/wAL6ujLMNt9sDshgLCLw9alVEP218ZVNL1bPtfbExZ/Qr
GuY3EJDLoICum6QnloPb8zJP7t35URPP2ql9ys/rNxz1eZ/DPqx/I6k0Fd5sny/W0xAdwInRymwg
cjq74aQUlkOROWv1HRdrmEE0ewHqRLEUAzkk0aKSULFI+q4PLKskH1LXjkUhRnjibQHb6RNTZSrs
sxr/rj6R3goqW/3sXjeXWenjUeNCBGF0gyjQiFaXtAX3y6LE6GAxjOywLf55PU9ONamco07EUZMg
KJNzYRMI0qwb0XdrfLxNWxp32lIXe1MqdfHf58kQtd2XyXBbB5DnubX1KWdWrWvqHNAZ6mmxUj8y
raN2npEKrN2N0GIqAEuGhxxhyaZRMX6D1DFB+JqXEPVbdKdz7csHNuChpZ0JQeSFdvz9NPyfzBK1
CwVLu2TFvKojuksO7eWgKitFeMFdq+w6UkVwN6XyKjF0ZPidlujiLSe/dJgVJTNmQFwuASfp+1aa
l7sPsXGGuUMfAkybrHHVsJSeU9Iqilg80VJ/Qp0A4385AX0goOSxdMFASxCupRFbIgAdBx/bflGr
EXoikcZ4zouvzqRHhysGp10oWL8YFuaPh43KHbn0wJK8i7XGnbFkcg4q4Nm7gXsrfm8c83jSVhEe
xA4TMfrVHFrcaR71dhObon1q4DLFv17hMgQnrcQjkTXAdkNCaf/y7PW9Dfnbsfkur29l43KaXrRg
fCMTdTqCjMU1wkSjztu6+ObqqRNmytaqtVdOvtoSere5CX4YtnQT7zxWNgsrPNpKtHeLflg3Ln1q
2kxAs7Rgfkqk989Fy5nGYLfaa1mT7VE+qCtVlRq6ke1Dfy7FrVg7u752bl5JyfgA9cOcn8r8YZHk
0x5HcS2VGl1KwPdvHeRVB7rpbDpzUzFGmBtivzR8NNByE8tMdOrdHfJJGozfXR3oFZ+UVMehqzVq
7r/bKYeNKaSMVqamXQAbJCrkK/MayU/QvhcEWSvcAJ7Gzp7v2DhkkOCROVNds0ccsz+Fvv1Em0xk
j//GWkS1OHJWjCKYfhijLFNFAIg91CBXP8VJRUk2aYT6ZzqhL3q+JIB5Ha8RUSytwHrdO23ch95b
8j4WKSsAkYs9cx4C0MZshkcPPrQwYkLn+aCSXBFD1YlC6wY+FFfsmLJi8Z9b+NTa2UxJqIqCCLD9
AuiS5h6khnt930DQ5dAb6fpzo7Vkt6L0AnVGGvhuF1BG8O6qikI6vQ8SeU3yw+VSBIap/cl4xgB/
VY+3f7vfqSUfkRwsZn18/SeUcIji7SiUuZ/JaHGoRUYRWKYV7IUJh3/mZVTNr1BOiFt3XPboKtry
tx3+bhN/Rv8Xi35LThbQu+Y+o92UGLOQyYj5rrO8iQUzHlrpXca7PGJFPf7QZdbJpNRvuIGPQLUB
32JRL183+9r21UyeKyCMcgCJ/hFUXOPfR3Ekc6dvBsMFASWO6SG6dcOnMoyi2+UYZ7VKRHX93Q9D
tvSVQELySs9C/EVVYvgWDCVNcSO+Bud19czV/N45P+jFTIUs6JN/YN1YdUmbWUdO3RCXG2tf5T3H
e61TxweAyPORQKkZJddiaWTeVwSsb99vMqM4fVotknC72vtWo1tbuQr0Gi8y9owNwERcYbA+qM6F
mNNSVTIMPzTyhAdTLT3SbK+dzWyn0y472mN9tVqzQPzXrFEwvlm7gt52jWmMPxcIFyvxwQGYJHd6
NntH+z/I8Xh4j5dmR9A0xhYpvZMv3QBnsGo0r8IKMkNpGdXIkIfL3+N/qHx87YbCblE5FsDclRlr
HIma1EdH15/gYdkQshLNrxsSMmUeYScjQip9ASsm5VLl4DsM5X1+2OTl7CRkANMLyxQdP4XhTwRL
Z0sZVUGP57Kx/0mE4wFBFH7BgOt0jydQPe8wXzsfj1zMwtG+LRuwZxBwmYDnexmOSuRZxximWmCS
O646dwa/ACzZ7GKciTR4x9IcKx8N91h5bN9d+CBXfl14rkPkTz7avZ7Nualele5pQccsYcvawXLv
YdUc1wDr7mSKRM5r8l6mEdpGkxQ/jM6TE0BbxZzI8xByzD6IbrkFLFBNa6U55rTNC053BN0w2KPv
xlRfuRT67x+P6YWoY/qJJVbvYfOq/q3R+VB5I7k+z423FgYNiSduvqoreeWmAPfKHICCmgYsTyvX
2aP4A7UfGBbOkjGPlySnZ/hfXgADD2RfmtdVa94M7UNOnNX517JspWp8fPDwCzXwgm0ZIZqfHbY2
++NkyBvEHJw2ZSxeT5CxaewQdtBoEFyDwkVXqVv+tHmEVXhssL8aLc0ell/ob30mPyLcVD+CkG1j
EAyydd8PPX3Hj3lTU2KB6lnbtIPZ3fkAYi+RBWYUUCdI9AoCiJ6F3Rs5okfqtICpk9wp+7hGrR0L
1YXMF+/wg9ntlkZtOdCC5EshOGMwuc4FdAIIdYWctqggBn+OVsAblAG0P3XEdrdnvLSzVCmf4m4z
YMfzkW9rm7BqDJ/iZw9g4cEGZ0ev5nhd7SnCEF3G1JSixvEJUkjLMasWWJ40gZ8CnkdeyYDFVJWz
WsI9f9m9EM7xvu1QN8TzJBD3PtIkA+cg4aN3Q0TWMUhLMnNB+RCQyzEeC5uWZVb0IpYsYHyuPF21
QYkrej0bFIqAyDdxtXMFThDrtaqiJu+RasGE7fxVtPa2ZR+n3zFcu5wfh/WqWHg3trPhKNs/8qMW
8wkkvB+gEH1Ivf62GiMrRfl3cft874eiWF2UyUl0Cg0N0o+ZM9yWs+V3ID1VW9vTU62kycgKtfiD
u9qxe62yyVVYxCDgWh+0nwT96IuNlMCOCJGSeNamuDekZzPTdlubGitjkEmI8+KF/L/tPXMdCpYQ
045sOmaOdQ0P0M6vRgPRE1KvNeygc0shnZb0YqjO6xHkwrxeE63opE/ZYYC7kOoL6wHJgBAc/F9+
7/B9BC9O89YlbUycVCvGxgUrRcbsYnMJCmws31aJNVVyWgdix1AFXakUcJ5K2roBytaXG9tA96UH
4PVhN9ZwF4JbD5XlBe0p4CaZ3pxT03oQyDQW2+wTHX4IuIULlCGzo+wOvt97Vil9IA/BEOF95GUr
kY3NamxSjA93CeS4ljflxWSr4vqknug99DpKco/i91/6+7DncDFtmqxSz7FIb2r2gxVsfKd7GdCc
fb8Zg5m5jJdc8ID1BCxN8ctNXnUlVcl1N2akymMm5B3tK3krGxR75y8Er5Mo1cZ7CnI96+9MRjUL
y6fcpedjkOk7NuumcWp69X9WIfznGesQ3Mno+GM7jG93cAlvnTAGvkgxaBhAjaP0zmPhwPRtGrXs
ImZx098YEr2vhx2ipkaLN1jDuf5xWPKJdV7ALiElURGxKcZ+H9DAr19W9bFEBuxtyZBlds0lSvME
NKZZHnyKW0IztpZAucM6HPTASZUfQWql8Msk/Q0loOO3Tu4UQ4cDWuQvJEdp48eOyRZG0QG94hyv
NTqe6lRzohzJcUBgb6oYgzbSi5ebPNbgRktDJsLA4DysXvWN30RBKXwuI8q9wbBAW6SOnjodJntV
JDcXHb4LB/WSxIJDOfXe9bzyXlgkCkjdqaYUG9rY0zRhxLXNbNa1ThezmrJP+XoXsmt0MCkyaOFb
lqqxueMAvQqTRI1UKceTnpMWxcl5jZdqJ4LzwYBtV4Y45IHYTgx7UFn3IWSWrj2o2qZHDQ3xkeHj
Bc1kSQ8TGNZTDEszu5Rl3phRll5bhTmAHZg2LJADqpJXuRr/an4JWqhwrRLbOs1EOLjrrGjfkYOe
YNXC5nDAKzHctvWLrLLnmEscLGL5DtGa0cgTLtboHbVpaOW5q8xL8FskZWoW8w1N5KQLMq2VWZAR
msa2rBDkBJjvocCyxCbvEidn0S8dDUXvJLFQNiuTxQPgP2M+4ncf4dM24tK3DBJoAUsj5jAe/adu
FwAIo8p+HiujvsGY2Xw9mThtb5uR/HqVxUY2+1Z6mQbqP91zKT84bzlQnozJLZ06L0m0/XusCXZ1
ZZ8+O/DVaf89mOT10+S6KHWRBJ0yi5ZhuzAIm2nvWbKS9fq9CcTsNW/NFMq24D9cGNBQhok7xMum
b4eQseDb3LDkNYzC6uEiBEZ4Ss83iZtGQswiDB4/YlAuTS9fJqbiRb6fmq4dzrz4g6NbNfhzDbYW
EzcSn1ZZJzmvsECLPVyYIab6GyOse5+jmbOODj1/bS8rWIyiFCenfPCz2G7Xp26gdRO9PcoMdM7l
QI3+xz5orOYOoUcAZ35Y1Hftf4tdOs8edUkaXcKBlj/jHhkk+bH4AO3PdEUCaf+UpA85viwGdOFO
2dh0aauEDVSu16z+3T+T47PBuj4YDA5tD4AJPLjKrYKtxODyFdE25oPBbvFhnOeH1FafWkt3lOwS
fAq7AupuUW4G3hqSa2lapLHCsOVImXYIGAMBsT3nUscJqxyjQBXEFQXPAdfIXBSs/LdGSDnGKWgn
qYEMG+9KdXFMvdyZBo0kPjAk8btaevwI+BfrJwhDTkM4m1GYyF8T1JqRzd15WDMTCCJX4kt691fS
xetScft+0qZenYGpQKb7oXC3n/4l/rxDGghM6YrtNJBi4rLjs9WZLt5oA5t5LdbTweR8D4AqOb/H
9RoGcmj4HCovKP8+olBbNpCYQJhWQCotd2BmX7nfMjKqQqBYXKUXSzTBPQDbPBlsaiaZTjYOIHPh
rvnZdC5G1MMsq2fScuU/LXOPuWz0uKPMHyXwyDWLpV8Cc1qZpUv811NnxzXXeK0cTLGGnSQyKnYA
6zaj+1+tBBUPmXTqkjkx8GWN5sFsZxyblCfdImCWjgfZjiZuAbrXRJaF4HYz/b85L1LvT/h98+ov
fGGSyxCGR+TOm7EIZdVB+wBxUz8ufIbhXLndgBSx3f7JyUIguJ1dsXjXw1OfeIra9GzPm5sPs2j3
eW3euD1W2tosYE0cKjJrwMkO1uC4Llv1+TJSMRr+ZcuP1CpfsrXnqBmiAIb+i8v2TeXorMGpyrW/
P5Y9lXxDXjmqg9UfAFJOqZbEjlH/AM3jpAJcv+5WS56ko59cb3py+ENhwRCJmyNHi04yFXFrrXyJ
m9bj35m9a4QPr7jkxO4y3BHgTUZFozy74motAoqvJZsR64J/04i9eYiaGzMORwug9mjOdvvYFecw
AdgpLO5JK73krpX1Z/uJfOwl5W+nbOKkwqKCy7i8bMVFZK8ga9h2NkS1f7p4yLa9Ekh07nbrOlHC
6KNMUiaEzSW5vQf4mO9KYYjql1OCcFn/EpIVWkhkF7y1qCYMsbRqb62yK7xGFab9z35EzF5vh2w2
qMr90LphDd1CJTiR/s57vy2vbDJVlAJcbuL98kUbf2ngqZlQW+fYnwem1IfcIK2qs8wKuUEqJQLj
haJlP5Y4uvFgkfu9oCXCC7Y1m3DjzKlY32DnLv+3oFpq1398FxqQ33771UoGjiSEu+YiOWwzpCB4
4JSe9e+6KuyR63ZnQhRcxYhJg9W3Dct9zZB06VYtJWmYWZ5U+rEZEXC/JRsfR819pVWH6TC5Cvyl
Ko+uNtYoPK2crcmF50AoWLi6XmqYwN9trLRrpWre+qN5lnrwzPJ774l/h57Rh8zBHXsjGYXl8nNy
pLan5/W88DEgmyFt2zsZsvdeeRk4i654p+7utal+0b0mB2OMOrT7l2sENAk07b/MTGCAmNjn74OR
vTfse0nyn+ICvG6Szu9VQxHpIYogICOOVR2Lrods22fl9cefqhmiDmFmuBx2lP/fHngVbKbpGiCn
FRE+vfSy+q3ukTH9aq7LrhWJXYanQ1D5D7IvnTE3q/+/nFErZR8Pz8Q2UNNhnoesvgPi2wOzyqmk
/ecIQdm2ylLZ4BhgaHXcbgSKvoaMLf9nkSJZPHPCc4nn6fXt/kvkiIatJ1ukmNr2BSjKR7kVIXeV
hHIv2gJ2l0+wypzGfyDbVy6WoozRr6ppOia/WnNsHXQuMbQporIVLS+Tcx66yL7BcUpmNZ7V85as
v2/uOkKnDjUStIJQsYRU61cjkfyRM8BW/IQwp/yezbj1XGATz2LgpLNEssTI1DiSZrB6OfLyZkwY
QsKd/nG6gwldRqhZ+AbbZ5cZVz3ldzqCrc2xEvJDotLADTrrR3sCJXaJIgpVgq2VJhiOqXmHnT2K
OVaoAUGVdd2AXsdOHtXQQk2pK4SkFmpUJm8AH690VDcM06BrQTiLb3h6QwPFLVBk7znuw7/mBq82
ALHamC2cO1FGIPHnsGeFXoZK3M/sCErQLVu9SNyit5phLPXcpvtC+M3jn/q9qXel2wEvxSJ0si+Q
I4JVS6R8mGmQXJ8eh966mzJ/+Q736Eg3lvuWRDD1OZvhE0oyop3SdZWkZ9Ctjrnfey/umFp7X9mo
bSDzfctLrfOr8eVE3+EjHhQwgObi6zCOuVEf31IAkfi7XVy3tR3MiJ12ndH5GNRy6x+toZw/E1k8
JUWdObppKPzljFHtaZCMjIBNQKOvz6Ur44PjmxYsNwZF7VnRyA+n4x5mpivR+vPOclu9Uh+XrbGL
m9/rF/AOvG8zB5+hrFBES2fIYrJSuXNriRDeMuyeytqqbux/AFOyzcSvB/iGztzZhZTp4UuthpWS
FvtgkdMaZxTWdItn5is9TaUdaou7+w5XsywGKRMOogpu9ywID4h/Nhze5x1fTYII5KUPJUIhrblt
z98bqP9D3yQyBbqkhrHCN9LSKkSN03uAAUoMyqk4ffiMnP7IDu62vWBkoQkwhnkjuA58tlWsbBNL
Lag/1XsS4nLQhC9WfQyhAN1IsWGQcn3LphGY4TXmPFypqFwDdPt0b4yvE5fHlaK5+G83vG6FP+5/
DCuikXh5B1tfb+8i3xK3rwY4r379TA3DDYflJXTUSm9rfFFuxdt6SOqogzTEJ+TjbixFIbS+qU7J
NrwJdCiakXEhht9AjR/gyNkGc/hl80IQ76HKOKtqTrDm8yJePj4m5zFDtRxWsMv7ieqv8iRjFKAI
K3GBFN951wmHICRdi5P+wMLHqkXNy+tzOXeNcgg4s2r12N1IgifNX/H8cELkyb3dnayXgsUYOqTI
oc0UAWM6CpE6lpemVvEYjDh21tOR8gucrJyHFN6MB2zN6hkAuxNSuwrz6LKQhPd6YCY+VH1nUKJA
p1uIPfncpjm1W7FyU1g7thgCHR+6U+IUmlnX9Igf8zwOj9DXt+t/N0H+J5vEms8kiRCiLIzZuVHw
0VAn/p3L/OaCsLA6jjpmo2wAMqiioJp3N5OY4LNGxp7JdWbwkO3asZJtPTD7LgAn+lJQLOrH5R5i
OT1aNa17u5R5eNlUC2SBIjkf3W224Xq6GDTT6RgNvWboFQe45mKJ9edd9sgL1YVSS11aWT3BSrv+
ye68x/5eQvkQpC4U8HTecXq/Gx3oNRWSfshxmPZB+aAUCd7pINiEqju7m2elx4QdkIZPw8bte2l3
NkFrZ79oKVgdw1nyW7boNb/7R8LyY7yzI0COA5qT9n3X+CxeN9VktoS2+uaEXeX4KnZe0I8WWlfs
XwfIg2npoS7ZjuHreVuYTsqCF29SlDo5hQTB5jobeGDl2eSOGxaFgb0x2veL1C5WgFVKCJWtYSAw
yDajeJpQNJvSHd/QPWdHRfbJ4/ZTkHvMX7cIumPHuIVemPBV3fe7idlz1n5lQDEV7x5C8zkT2d3s
3IzNmCrvwPyH0LvMwmQiZ41OdjjqLYW/ru9tl/XuoxaH2rABGReRzy+fGwz5iL/P5P+xmQT8RTi1
GCMVtcexT0XKXzwFabNWmHIkL0S+zvLlthxMkAo5R6sAsRqo6YpTWv0zKT0cRMv9CWAo8EGvt6nW
d5cYzCrax4pIwhVJX+sD6+HbbzxEibpH6w05i6tEo6+1dtDFaRV6qxLhTd3VUAB1f4bdnZu6kWjs
qsdlSwTCdVdwcA2iXPx0DFRJHwUQ5VtJ0k81x1sylZgt3xScSElbEAk6WYpYKdwjciKGWOVt6FvK
lfG/XuyTeplP4wxheZ1KB+ni82EyOVP1wqn7dQXQuKIqYIKC97IgS1uCvB7If5PodmfoPOlT5OQm
wCAH+ms248U7GCesQrtLjhV/hcjmjx0NGzJPr6FT/512TiJo32HdsK/eUHNSagtpBFYwA1v0pord
UXfyYG2DDp6lzY34LgbKws0rarjuDLTVxL6kFjtlaQqjqTXLwUyFk8LZ6X3GPqfl15SCx+5+jkBb
lXqd+g7TGFBBG0YVa6dc4N81YRY0RpehcMR2MHgpfmPKRraUIhrvBR3zZhr8TrQI2xily2BlUvle
ivvUG76EpJJwC0ndbyuMPu/C6XxPQ54rt5cRyWfTqPKKO7nglAOZ2xUfyG0Wwd46+hmUoxdCcrOc
v3TfNPBr0LyguvobsGxY8xOT7b2rcPeF7aLFVAhABgsK+L+j9mbGw7yICqOYtf7ULM+HlMvikfkd
Lqf/tqiXIzNBsu0ucPg9Qe/mQhrgva0iV96rMown9tb5aeXsWiJnydA/5AReSkK4meReCsB0kEqi
PQGeo41lS9JB3tOjXovuNODllCSgMQydI8lXjgdfiSJf4hrgutGT/9MYBQVt5jQvav3iRvOLBmwN
au7NlF462pRzubMZ/affc3sIRTFWBfwnsFnAO0nRGQF2YteN5Q2PqfI5hL6HQ4PWPx6wfAOJ1ODV
FIzQ+zvkiZao/yjvwAoIRHiyVVmygWAPWXzuliYiRCrJFphd4vEe0eels9smCCaca+8Np+LP7U0h
Eg6jzs8prjyURYdmb5FUj30/hwTw4jYC8pqRjGDYUlKkKjNddHUMcaVtQfAdFr4CyG4vPJQuBviD
MQf2lrb0gKlM4pPejPOPTwDSnemJhXxFE4O/rd4MsvzcSwfrS/RX8RMi8gkeJI2fsXo8CvwjTnDr
GnDqL95XyrlKNT5tYO8guEmzsyLdGmEjGzmQQQu5s2W5ZiMBotCRFiMJ1I44gzu5+VuNJXmg+o6Q
0mOkuSYojc/7/NWM8HuhlIMwrlrkkHCcekU5B+xh/xcUK28Ua+sexFI03xM2lUYxWs5w7RjQzLGi
JIIK3MLoiBSfJS3D/7f0YkS4PI+PyOrXNx7isfbZZBFU2YjbTvtgUc6Wd2oeZo94ym4QsKLfeujX
7lXM9bwppmhtqXpl/Ec3a6CqgmxpXKApqCNPcZsSTSM7yOmDatPuhvn4t4Q4MguvlvUM5r9LPhKt
p8SmHjrUIpBevG+kyiMTLYHFmEm0PXsRq9wchAjraUmxWYaZYZMeMSNRBjZJdv8HEkJeZb4GiFdy
hzqXosoUn9NcKnn7oWlPAMMTMt1YlT8aiSTXbf0xvnO+bjuSck0uQOQpV0vSQ0nvQwnASNz5B0aD
EubMVbdUzBXag0tbR+ER1Bv/aPwAq12ZX4aL7eRcwPBZMN22crmsdvRzDYWJCJjd9W/2/szqaLoC
w9ndvjs9YuCXYJ15EM0WdQrFnWwKYApWyGbFo103PVet+QUdShFn6DQQmzjiUHM/cEDyO6D+hEYc
3Dc8265UJjpIsy6h/mXMQTe6n6Z5F++IB8nz0kKDN974bpFzSu7AwXr04w/VBv4AmxJGP8cX6qNw
mQLupO2ZZZNjLI1f85ZXoQu9a4dwBkZJI3HhIe4JUKNgxZ+IPtT9UpolQSW+eQ/Gj6F9lb6sztC0
IixLOwqaZI0YEwN9LTa3o80PLUEvEfgcnndQXyjiaeHSkLDlP4I74UMPhX9Lc7Mnq+wIAX7sBq5y
2IcMCztMWqvj7Q1b/MSOQtA06jK5xcbOo+a3p/msQk6vN8DaJCcPg5upQ1Wn2CSYNTIwY64bA2cd
QpuMGG7sH3j92oSdAQtKGvrxo4nAgdWrf/gRDuPKAIPsRgGZXdKhdLl40a5y8xCxTEtva3/x3PiR
pQXwcOqBeUJ/WB/dToxT8W5sLZ9K3Yy8vEI05dH7Vqf7MIg+U8SakSwLcHoFYDt5ceMiu+GOzRhh
eFYE5gdPRJj7VSvlnBs/WfmytbRiUvZ7JRJNrqyqdAW5C0u1kaHgtCuwod71X529gCDwVKHQianL
l/g1PB4C+TMicu2dPdEO0NONaWAhZ4WQTYlsxZTpJfM4C/Vf7Om4rcklLGQF2dZxp4qCGDJqEatv
PA0SjO/winfYKMvlIUDusgFj9bzMjz8Ot1PvAE2Vf1W2tH+QNKKhoNW6kXX54EB2CbsHDcLXupwQ
e06IXd1oYiBpSh1QghbrMZxYF7rA5xTnnh17iKVPXJtQI6G73VhZiy1lB2PCHu+P6jZzAMd4Pr3a
kYIhY+sVUinFoiVJVLBQ7S6ERuLIEoFj884MIOddESTkhq+ZgM6TZpbO+Yc79F2ocYosf+mzoJyt
YEOMi+IzsZ/sLRRUUBgWPjTvr91QDMvli813M5gKS68DfsNgvxt5/zS82WywmNMqaeWkvmBEBEwH
Ri4g9AmMH01VN2EDMEMYDx79MgiXxudXiw3msybmTRts0VhbIbcLDEc9k2msjS83MEwjAl7mYE8i
Qxx3SnzFyTGzX9+XSy7f4+dI64VJ4NURnsnPJMGUWYoK/vfcznlKQ+Sk6n5KUHloO62DJfswOscG
ASIc3ZAk17uUcPGKiy63zkQMbSdz+qx8pNnb6nqPILOQWAiqNPC0eFsdA+Mm+PCpkBO4Ql3CDrL2
V3/zVbnCmiFgqQ3d82CLssYdNWxSylCv+rjpdnCa+mOo839TXdppdthM7kkP8G5yNu2OzseWpkCA
nDt1MXxr9AjzxlETV5zBxkPee1do13k3uz80XnRRQEmJH6u6yVWPfhx86Mo9UHJMr/zOgdUd65/b
J0LM1RdOvaumaf3+a/4LPxsSuSyv1Q9wYwK/C70R9LTG2kdqrGFtS7w1rOrerRaVbzjqqGCW0DWG
2CasgrhBt+P9Z6q9UfsPqV7O5Sr0Rssg3rbkjsy8bAwyDDCynVfAfy2lGaTW6FlKpi+hKj/hiOC0
hn9Pdc8JICyojWLtdlphW81cjmk8494E0MrKiS2g7cNwTyRJuVmpH/a4qJqrQ6C+AlahUu0D8ISy
O3Ba8Sq+JdLMp7mUOfuCbgmeRM8yT0jg8PoguMAllHCEUiH+HrrSelo/kRy+AYFd48Nvkqg5hu+q
rY7FiJpIOUKc0FmLwvuTlob0UVE9OcKsOUqXJP4/bD/3KTbBZEZaynnI9h87b0MYX7g1ZrLdfCMn
XdavLXWWCOQH2TifUBMRd+ClA08IZp1KFztkgQpfZZqeOplQvHGqImLYNGlBEuUzqrpRocjbITuZ
lrAg4ZmndT4K6ElgUcUYU/mhVmasu7N+gL2zIjp2E4u+0U1w/JsaoXmVqPaeWb7V3s39A/s72h+a
Yo92Kp3F7qCpbw7lSr7M5tEKeiKC7QdsiF1ifvNcU7bZGYZenLHaZlo9e46GiNSr2bTA/a1RTrPe
H2SXn8m5Np2o6Rio569Y/6p6OKk093SyT2Dwwzy3n8yQXXbof+fE7rAq8O0WPPelqb0rA0thtqtt
qVSD8RKF4Z0jsIvsQmM7Dtd98Vk/fzFgaNIMSKWnpdv63HLeLBptmH7TydktkYPUCX1P/YaBYX5L
vsC/WGVv+JofZV8s3Fp/oSMHwe/G6/oOAUcATa4lUz3Z0xPTMyQU8MQ6Znz1xrpjeZIx6DRKP8wN
qQR6Z0fZeMutUmhbXsfegq1WwpAxF63JM0IoE9JtUxxyd7KPUBNV99HSKBAtu11BcoPZQdXiPz5O
CZRmycjx1OG2oo2s78dZAzKbAozRQE2ilLRwB3ygtxTDln6KASH6bbeAdoCjo9TUcDN8ECBzGa+M
nPlBKmIBlAmlDGGkotX+qDkux0jzI8r6e6R1p+2ZsDSvg9E1u1SedroauFPwWSnVq11E3HdaDGMx
C0bMsDqTM0I1CNwvxLEH8lxvOObcJV9kHkhbwJXgZUqXnLumLU6YvQqaIHw4EqNiotCBGg/qXjOr
7kEVaqt0JM3eL1bVb/Fh16oqKT9zkgEVpV7dc1tL+4wkjOvWxWiN4UBTaCoQpwIS9O5r5AXKgb8B
gF6GDVmXRgtjN2PqMQ3v80pmgk49FjFNYwPb8hcLpFgDWYSKWXKP0t3Tp4So60uEYbnkysoLf+k/
1IggKkKiYKpADexldGGB9k/TjQPIshGkWJD87sqsVEZJpxvLED9WanAvz7qWUFK0aXcXqgE5OSqT
wh4NQrgsNVtvSFKaNYoUnQGFtlpJjxIt+lAOepSxY3A1odIfokIEoVV6yW6ZUHScuYbHjYYSsPqh
9BmpcC4t/5fwmVF8o0RiSnudwS3dP5jWdIzr7TT+AbQYlcOcptREX0n0GgeDosabWdx4QV0gLEks
EAzwZmri8/SWrmoT4I/53DMq7eyR47jk3btzeBsuPw0IOQ110bMyArNKCR+9kPEocuY2yND0enVM
KSubNCOciRLN0uaHy9fxnrAwAZi6SI3chvBE14lbPyiJYQl10W1L61CUPz0Le0qfdTM6XIC6paM8
K8EmMSlmvKWnJReX1GZmePuAguXxNc20Hj84L4ba3JDJ39+MF7BKYhuFwUaAnEWMKAk803E60DvF
g+RN43iNqw5kWLX3HOThg2cj0YD7fSLOkj5aoKaovtO20ZxxsxdPPRU7ia4X878gFctYw/Pr4sOA
oqebttXW1MqAwrXKc7945aU1b63Jn7LYwU+fnYSy4akvI+csn2i010aDDQuiRwvuTnDxckUB8dKG
QIzHndBcOuTpmS+Mgjj+t+nW8YZxUC28yPkHdkTcTd+x3hRPcW7ZNa52t8wcWxYcfkJZlN21i4YI
D20kpuWqmI81x4oNiWQVRlIzDsVu1z0Kt/PaAf9ZJZi7rtKxCJfRrJ/nKwgMpFo49k/os9K58Ja0
3/G9KUY/Hvi5AyPMelREB2aeqf9mqAcrwa+Ys0uQt5mrXo95+31j4kHGE+nNNATgOTJyUbiubCgr
zGANILK9IbjVrZ+fQWI6Otzab0uDy5KRYVpzuDqCo86msiIj+/5zbbcuZPE1vhp+gw8QENauFHSK
eGfSB69Web9zBe2I3wUAkSUzRMmgQFrFWyWbV/9HAQVi9Y0SFEw1laMM3CHKjBdikr43ygty51Kj
PH1rU91n1ajgFuJycDedbLYFvtj9k6DcMnVvfoj6YHpxHd9tg9zBHCwxkc8uF5cxjbOW5hO5YPEu
P0fD5Brg3TMmy9dOo96i7zlgbZmt0vRlAeLJOkZiUCDwKh8rXgGk+db1lHCOZW6yOiz2T4Dou9YJ
y8akFxjmZpPnibdr5FldWUQKGLq0fHrrtaRh0UM9r3CG4CRwevj5V85+a/f5urOZhLKW2rkvQyEs
0QY4/rC60ZOsYGlrK/fXgJ+CUb+yf4cRYFMmupszXlIOUqEYVysievwX39wVuhBHZ7TK4iwhhF7r
0FqfX9tXykanZ/JJ7EWrrThYykranswe8FELRvJ965wVBeplXdk1MmqnOn9bsxNpLGe62wfyDb41
s5mi56Oj6MhVAw2zHde8kA0SMVV49VWddwJVQl5ZXYT+xVsZ8AhvHEDIHazFSM50ml1xPY7fXuVW
7bKmDuuxvue6pK//6uZMrzcM2evrPtf5sTLBSKTFQBhy9NsV9vEqp6JzZoXu1ixy5tmBirdCFZYz
4iM+VRNiogfedFExI0SZgnyYend+g0eHD6LidWwEp/3YMeNDNTVcerAL5CeihAv3F/KdwQ7hTAH1
5zgkzMiU/c8JxtZ0NotRjc8v4ew1FXCFEIeQgmm30D2ZeMjAPRnIPWAME35WcHb+PYJUxX/e1P7V
9IjgA2qozmylR7eO/NhIaMMFIILX1SaDbf9AC3K7Ro/PGnmVEHTGDT0VVLgR2OaDixZC5YwTBqfr
+GgZaJGZ3ZdM4vgbWjR0/WX3XSc/xgXxZlGcx59SDHX3qTFuoDEEECjA6HUiSYT5iH+hn+cI57w6
//gpdF8DPAkYfIEDNAd9d9QrHs5uBIk1RTpqVpA2lQ1rqEX6B7+q6aexYew1210h2ZqgyNpEl0Vx
hJg5ExCVdTrKDUt91knHF6l30yjqwlTGqH6HZ5+QN4owh/QGR0YvRM9JpmjUKfT3edFr+wKGqVwb
hAMOk6E8Ykmov1TDe8WDjNxuhRIMrGK2whzm8I5U5PYGvXHy2IUmktuluKzINajEqMGshAEg37Lb
vps7+5VYmJlKvSUR0sCUJKkCfAG9bDUWyijmsbXGPDt9uTFx+XNugouIPZkx9p8QidmylJnL9IWG
8TgcVtLewdmIQumYkftxsmViTWkNsJ1ypeNaTmtLy51wo6F2q6cbLRBkHmbUgja9cO+bKpl/pcr0
c/lb96pLrcdmVoFr5Sxugr1rtZ2+NVnxC9NaYRkQFmtpSEsroYCzbDvAuPAOYpC/OQRxyXR9TFGI
FHniWSEjfMzXYrfBhYZwtOpChGduohZi7mM1JroZKqyNXKtAv7AiLh9MakeuiWbMEz4gnLhjjZiY
DWXAb4Wjyx+MFb7oFsFeyWGR8Ny7l+d48xVMvVzSUyme0iGNhbO9QZDl14WSrhSfN9DAmbTnSF5e
LiN3rEVOU9+RRF2gm0N5aEOZ7PH5QJuayK0NtwugPwHmCzxEPqvoWl/dfU612vv7fFK+xybunv6y
DwA4oYwXdogJd2IIVMSK9iLy3t5mI79X5QOaNCvfWBrGitYOwOIL/3dt4yax0WPmFTThAWcegagR
mMWjRJLz4lu66A3xkW/wBwKcRIWezPZBNhZG1QYI5Zb57OByvj7Q1EZ7oCkn1S5GHMOY5bK85XOh
Qtf4iNqNLj7XMIymXlelhllVIILrQi9unw68BAsLks8H5HP9oLumB+XnlFAaphoQT8U7Ks2EJaAw
q8lZ2di6a7aYFkXHaqwvv6VCXfpOmZPypRwxUIFYQztwUsPaEfyl9IqSffPpL4SwO3KKMMVi1tIZ
H74iNr50EKrMlq3Q0Un1pCy0LDdSbux9w86iqD9sk55RAqwYBM3PGUQ5SbLJbDGQoo1umbyQbSXi
NIg3ThzQgDKr6S458TknOFVOecOPm9+MMqC8dJf+8HradWvX42g5pBLVUc/m0Sxvi35/eQi7ZZWy
+NAGXYMsvsWVlKGUofWLf8MZsoxz4+KT6VVlRllBnwB3bWf1mocIdLHmqL+ev84rRntLlgfwTBuv
aV8pFyL4QMftX7FB8AKQ3NHEZSWxLwNpuyS5/twcQtp6m1Z/uQ/b5Fgg+9jq3Jj6LqI3JnBb8VOq
HefMSznqOoGoeyj0wc9g+4QGN0an7Eo7kbvVGFDpM9ol+TXE3zsQ0AuLR82iNm/HZZDyu1QPz327
1Ec9gCshLx3WnURGIf9qC6rF4hqlUllnrwnPRDw/LNAaGmzVeO2llcmfGhSXULn6+EkrPWFybz2i
Ka3Uu0zw4bYHVwMN46SJj2iytibS8BG1Fz3su+oECcnochmDZBhFJ3w/E9lV/r5wMl9I8ttV8KW+
wELXQKX8/flWM0cN9eBiBeyi/u/q+spaQZpoNh1OWoOCGUVvXBfMLrVlZZA4axdoNy5o7d/W/12V
fuIzMgtYBhNHpstdh2jv6wPeaf/7kXbxapZ/cr6WvMRhrgs6D9RE1JQcQ9vCBeWXGR+OCXjyCoAY
BPfCY/9q/D2rV00S2BL9VQr3CjNW872qlFfC8QJDUncaGy6JlkUn0UM/NB1HL3F4bnI8ASCXJmy9
+0mJAmAvoJVgng+SgEtudZ9TJUmVE+nTn1mSTj3ZO9FclDcHjFGb0vVCAtGCo6AN6CUvMur0cUq+
5Bljkki2As8D2wfBLd2HhcKMMxQBhNDuESsO1QO4ZNo6fydaBT3wrygfJPQQ3O4xSCB2crfz32Tq
uSvRkIzk/44c9BvFq0njYp6KcvcWok5/F3Ts2VEVvCCinYVdM/NL+IYQLAgiX03Z2INgoRKpvvAs
brHvzu9rmsHwGHSP8mxZTNQCyqNgSu/sNqShtEtQtLTzhkDdiUos6qpAwihQfajyu1bj851A9o+5
pOzbhft1mTFf79CCJp8z0X4yTN7x1FHQxBNAh79Oz6zimDbWMEGQ0ZS9HHATqY2ey/2k7MSxIZqI
0AFF1LJRW0kUwlAKF70/1qnYk6WF13rkse46W9tw6Xy/e9qVPOvxmqgdhDO2Pq8m49z5HrRJg1Ry
C5tL6rL7Y2ZAoYJXWPU+8FCh3BgQlOWWBb3DXDRtuzWAmUc3BX7xHco5Nnsz7ml86tFT9Pg/p8KE
rrUKeto2Z2fMgMvCuu1C1UzqhRyzurxNze5y2Zhc2ms347RdOLWEw0VHAb6yuBTh5V3Cyb7PYhH1
/1JuaTm5ZVWGISotQXc9U2EsC4jynDxxfdTnWedcEpnc+YVQAXVxiyKkKtgNZeabQi1Bx+u7OmRg
9UvVacTjxB5E4ycDAzSe7ubRcupgMMBlaq7XkIwQwA3Hyzvn7UYQEYEbhILcdgLuxoaw0DYdUiH2
rKFxFljf1iGcMrTWUV+iQAZc/YXgOTlehbuMxsAuFKK+dTDReO+JXcy3nB1uz34tlQWFDfKv/7BI
u2A6B3aGSpx1nGmi9dauhoJE+qMbFzmTStOseebASadte0CE9ESUmjapNt5riQYKmSmZPT0EFvGp
LI/FTvGdn3PFciCHDIMgokBHjYRjQyoQgYkADIfg57Hv4hBsWO5HU8+eZEptqPD6HNBm4cT2n0/Q
CKD7VzagOmVFp98LfUyMYdQgRfj79VV5uKqhJwtS+shX6x9d/tAGRWmC5t5tI6HQZVntmPmlCaaj
0dsg/SOqGMRYX1VD5a8RxnVcB4o5Zrw76v/hMVCDm5In4XnFM0azAQTpWoLpW3xBUTmlK6Vng7m+
At6W3cf4F1T2j5ZOtR//vCXPZfkLShCkwN9QZsFvl/uBBDMQ/p3WQkPHFcxUJNE1JECPNK3U6zLy
eX56D7/+XRR3Asqwy1nFXlRJbTphVgxCTMnr0xCQGIK/BeCmWGXv5IaJcq0R9RW1faNh+5k+NHmg
i76H5E7iER80z8uGVQbxkvSkP8KkT1H4fyzyv1Xv+cPOMWuoq/G5TVB1wIK+VaMk4k3+izMPix9P
jKcwLdYJU9eK2Z+z4JXvPwqJzTvxZOtwZf5qqCS5FUYVB+PBOvRdbt51eSzBujP5/4O9qhID9mNx
mjj4sq1Zkgmre7EhqIXEJd/senEY2+DJ/c0tFdcukjCqi/94QcRd8y50cSuIzbF54DuXnkwBISQ8
9vqOwUIp0bCAbQPeBsDdiDfd8T0TLwlez9HenHo7Y3Ls24w9iX/dB94on5JclwkRKqhGHnU3mHgk
MxjV4b8Xe0bbs914je+o3v3hdvdm0VtVYye1vNRamoC9ywlGUp7+uN2BcU/x12Je8wfJuaE3rUhN
1RmPfCdoGKhsmBdJLorXUC+XpsD5i68VryFEQe2FF+gPMtmWE9tJNspb4wbl74gt2e3+FH0viQ8H
b3oahrJHE9vPqWU41pG4joG7qPESqLyJbO+a18x2La4WWAziMc0w4pi4npZ5PIimgq/EyrNCTbEu
xGXi8nBrE9AnOx2naZHyb5FwIEyuxrbIOr1kaSgMcPlygF1ZYUR27qdzd7dnIoUQKFUB0ujKLuOF
ztu6t9183CVZKdO4TFEFmkp/x4s9crCKw8RYNWsRliBd+soeVkFeo4s70LixlSGhojDW2y1PLvu5
lIcSS6I8bJt4rDWugiGt6ctRfcw2k5q3U/uXM4JAPgivEvCqqWhje03/5xLmDecXyUmlXHtod8Hv
yen2/Omn+6s9hXPo0NSHoQYhjsOPG77JC6c+vmkeGKK6wAMAws+m7TctkfV8TqJvhq0LnyCKmNjC
84K873qZ3E6aiYjdKLi3XPDdgaUGTINRh0dwQ0ocVnwtfDGm5M5nwANQUjRl9uxA5+Zaw3I1vk86
D3R/Cn+YoVh5WURwXskeoUgcQn5XEHSf3MS2Le4JoO6zIkCdNmshoAP6W4y9LVUw7Ap0irmagdS6
eMLQl58aa+6toNfUYbqELE2tNPsAhmKISQW18lTm6Zfsd+E3wxy69k/E9aebu3LNVaDPV4pNt2Jf
sQOzIIjYU0QMQbmRbT6ylR68OiE7zMNTcyjESjn9CvNNenUVaA2oZCyj7hRts0giFkXgxdNlPQ50
Jiz5jYkovOqBZmzGqBX1c2Fj4P/zpiTLgHOWAtph8QfTT0Wfosm3uk8R4cdjnzM72A4UjCtrRKwt
ZikPkAgKpWWRiv4B6pvC4DqiOPLwNACChYHZyEP9kYFXuqO5IdkAj7iy7eTnfIctir+J4dwXgjG8
6e2Nw1byGbuJ8iiKtfehCBGu6TGV1L7/Pu9H2mhrzKUWovVMFjT+MddFwQw9zhvFwku5BfVs+sIJ
z34EW0n9ncbrvf9N+RUZXPoqFrMZ9XAaDf8h2hHONyluqrueJAhXytyyfNaQ2bggeNmW7gXqnnfx
/VlvRrMW4QLeNPJPQiiBKd65G0uLrR9/YLraEn0yZVBYnEzlX20CKpkJQ3B4Q4NHhVyco+IMoY3B
jMMKy1bAYZQxQOSCaphBNqNaiFfqTFczLLW1qBpAMrEdZaIToeT9ksS+wUtAVJJA12A0Z0tE3AW9
QQvHXqLzbODz+jhj26p7qYKNQFO5HruCVBBJLVD6FxT4Qg1WQ70cVf5wYH5Nl56Xd9vG3YV/rio9
0lAGt0uEkOXhuKCvHHe3PpMDbniYvZw0cP5wjJWXI4evzh+zDDsu29QbeoEnGUfDEo+xLE9M33KX
3/Bg/wwQbqD7cZwQhRD/T5rVg88N38s6UYHOQqTOgy2B6y9k8swkEmyWnhlVxtrq5m43gtljobIf
E1qAhrWPeB+etedHIT4ruWvIyt3i4V1px5da7pM5XtF8gLBoXm3t0JVKiolwMvJ/QtMX+kKOe2rv
O7pqSKuUf2TpBFhrc0zQy4wvyNxq6/4DWyk8D55iRnu8N/urdbFOqLN6gW33s3icDRhWdcRp9Rsl
OwtBYXlVvQl+CJH5J9btCERQmarStodqcMOdA1sDrnUCDg1o6pDtGxjgetOWlUAELgMf4/k4jx6O
P5bh9iHxAQDPv9VYJzHIVDHucVBwExtCYVscBoZjpwIy/TiTZcW5Ob4ELdIgEAzQXZUwcQ69JoQ2
tpCM4FYOAE4+dNxTQYBL1WEngzCzTA66wR3G8SfH9YLm2c0miNhbHQZjCZl03WVpMB9YvJ1IXiYV
HEsiAbmiorY6OAFR46T567/yHRVAMQHRqtMfgy0XyPIZrmSRe8ow3TfRdbPuLsrOTZFf6JMYdZk9
IizmvUJ1haQoTDv2mxE8aZGdXdlXWvdGXRjt6SAHddic2/UmR4GNvgP2XAS5kspG2r6d7bXB625X
0uFvBJ3iXQh53zC/rO91K9a9zFXrO/hrk0GxNgDcXCU6ofbUWPm74zM8ffc3s6rbqq3+J4Cq7H3m
MrkO7EhRuiynUypIOixkRnpU4xpqkEqt/ySfg1k4CVE3hC1O+w+6MjMl4UUsBk3jj85seKU+HrgV
kG4Ig5p1h0vi4whrv7KxMPMyIHiIWBb1/p5c7k9ac1TZMZnlK+zd5IELdsLzRfz4GQ1ZdhbnjwFD
cH/QFGg1gxdnIdo+tq8DkNDliem76ZPgJX6DA347kcRuUexq9PP9muRmLN9r2sWiYJ3CU3LH6gIp
ZNtSRLlBkc1gukIAMzelNAmrou0wCGevGuhXAlrlXhDw7B7Fh0RWYs0fffuZjxAyHRx16CykIXxi
Qp1Lyz7SQ3CAT85y5LV9UPW05niw4WigpXLpn+cdtw2uwGl7v7PIxgSryDIk4Yzx3FEEMzd/J1+5
xr3HWfdkg3vEjlXKK8MUK84/GbyS7aHqJ9RVy6VbzCcJOG8mp+0i8d4ICA/f6+FuITBhatcOliqS
Ve//i7T/bAunQv80c6EwIX58Wo9cJnEl6ssvh1SEvayFkZZr1uNNePXvhccZn8ZFNsdPUZBCw40j
W3UEqn9HK6vuothgtn1rEtOcph8+NZC0plI1sXyoD2boNaxM8AjKYZruuGDx9L8ZbIT4ORs/gwMr
nvT8a3YPiICzOmdDgF0qUeHBAONBZSNrx37MVvkoJpiPh1W5zF8qzQZ9RJgOeVgJGwgu7/4HQmpd
1H6HuMITxwqv9zHdUam2b+hE8/fVlHsxFQAon+RtIbUYlw1BgDev0wQCZNWB/P0LW7BYQ6mGndqs
B2BAirBKAaYTRTyghljb+FCWNNyyiax0QcjdIFJAMTcbJw2QpM01s4I4k7z1SMniYZXZTIM/ynwA
8J1CvUCyDdhXGe0pzP0D95mTO1n4VQYAeoVCiJnklUs/w4c/6OAmpPonD3ytruMu047QdDB/hm5Y
J9zf6Z/+1IqX2/1iiP6q3mP+YHi35es/R9AoF6ccjXO7rMTofTrLDqHuaVzZqlRuA4yYZKKsSdYF
OGJKNWm/+ddePQ8nyzSnSQbVz723fIsjOQI8ngnq7gije+f5HadCm8cEV91Dl/AhpMNVcIze9Pfe
eqBrRiVrLJK9gJ9w8eftfnmhEAnA7AK2N+vB+ADbE9Zg7N7F8Hxa3NrNAAi0LewjD8O66k7ujsNZ
Sk4ilLjyGvhiDPaeUjhpaiPArpAnkZR5pbX8vN/SONctgHjjJJEhM33ogsgTVSR6ciKDhiA1997i
irks6nUtt6Xd53VB/0xli2aKHL5zGmeCTkl0Mn2E4/UUanGaR+feqNEtrY5Qaj6LC27HfIGX+dnb
4qYVEu/axvX1unR06UdDCW83UJoMck/JtV0gEw+GdZ17NoFiHb2SBm/VcWkyGLRX2Cdxk+F8bgwt
OfQkmHikBWKFXB0PVnfFqADTMHq+mPTUQvTzQeLhFA3IVwhmvHtRt5T5HkjLqhAnrovUFwJ+wNuW
Eo0tHHXGiI4gzRGux9Om1kz/gCr5N+GmBASi+dwcFAkG2rTGl+Qpxu+CBmEGh2CuDD1QoAKRD7qs
TIb6D1Qlm1XpDwPejZJmXCJaD0BnbUjVQneeB3F2vbvCmgUzKw/CiHyBLeqqZ+gRlfUxq2A4ulej
ASZsd+G5v/QDDRuOHOrFMXjn7Ufh2GRhRzU8LZrr9z20hAu6w57KYGTenRy4018qjpyyV69a7vl0
4TlIfHuEpTIlKo09HbcxpMooFcNtcrocH+w+jJ/fTL39ImyuvDXHChif3QIdPm9RFDTAr4S1GdVa
NQg9SF/N/e96AKs1o/EyUKzYBc7t9i/yrKInEsXypN+Zgpk6sCYZ59romdhasnz4flxm1B4Gm1CL
cMiWyY9MYNwgN88w4QQALZ5L1jBm+jBbZdIeA0XFOSqhTTbKr3LprUyULtCJeOFuZQK3kaAywAf0
dDhCbqrAQwMWStiqVrTjnpJzHMyhTRqqYQd5vrNJ09AxMcf6y25RpS1jLhlYnhnX3NDKYvDx7PlV
LEv9NLOewH0K6u/rtJYMnANUOeEVKEDhJrePE9PaDNwrTAz4LgQV+uA0dyk8wn1VzX8xdCQEOYhJ
Gjw2BhnvHdajgWVnBAiK47BTCP9sVLUf8kfBLpvZcRuoraGxHwJjXuSkHe33U0MqmNVM7j1Hyr97
GC0T6i9rAsIAzK8Jh0K7oLpzS4RABBW0tKYlf+LXyBYqbihbYWuRlNPmcUvbtP74qZFTcqC4ijzK
dDq7MNmZgPlYrXa1FVvzurT/XuBq27Xgco/5huv7f7x2U+iy00NppSsDxWUSW0nybIJw8YfNJMkD
LdfBGF0z1K//25Ut4SFKa8napb9OWR/uosbhTlxtMkoIC7aQVBkLL5oiv9R3QSlQoQX25YZ1gqo3
yVxu7CbxfPkK0oHySPw04bht9/zfBMkQDI6aswf3rajf/LJRfwjHFV5DE1edKYeUqPasSNTFvSNs
v+5to86cukxovo4oAZBApyg5uDHGbvtuwPcApFQoag1LDVcKFgOzummzq3A/nYVOSA+wT3GYyHyQ
Af1h40OMIB6Klxq0IMO8mDe75+OU0x0YjWX3EN7b/BcBJA3nkPcXRIhIpPMG6aPP5SQ5sUOLp5H3
FiYV+WI+Jt3Ic3oCJn/ajDGA893rh7ErHMc67IO+UTqSq8uve9pRIvm+Pj00Bo1OpYTw8uQN4NDu
LOLnrihTwV/RFliLrbZTRJLFXi/Ti8vNt4/QNgZ1WKQLkaRa2sAWgObsr/XLNgKkHYHkIosJx+dg
zbjcBD8mdAUQxdr2VepaSV3qwTpNsDH0wI6I6zkslbDG0zm0QBL9QNYrrjQdhAsyGMzx23AMCDga
kRhdqeWyL4krnCjJvCaKmOzS6rop2Jwjap0PdzjUJV39C0jVb/BKiaN7ucGl6ipeLP4Qw+5rGCco
SUeIwhWQh7v75AkACCZBnAR3+mjNjn3zII5QcTNj+jNWcsKMzXsrYiI0uMI2BxGV8Z/LeVOJ3rwt
JAF9dzgie0nHcCKRcIw8CDXMqPZidVzv5Bhjj8z2iS+wSw+TLSWBRiUUi7+eoJmn7OG/aJKCzojY
vGj0gYaO9to3wwOljXGzOzo+jtC3ZBEAVgYj2VLK8SMAh1QTCaWuChnRxHxNB3GKWDoi3aRsoX4u
f/lEMDv9Ddn8Wmk1T7PGmLz6wwnYUnJi63rqMA53IYjW5dKaKZpaWomy1aHqPWO7DREU4dz9R+/1
tlCNJ4vmeocfn3N/523OWuKjsSm+5V+Ax79Gw4XXTmu8QiUe7WJuZ3mTLe/TKdarxb/F7XVGDyGC
OL9zkH9z7b5Jo8GtGLu2WJhhH9blP/T+LB9vdKQR0jrxHQrBVYGlhLdeIIEml3CCVW3atmauFnhC
zaBt2+06cdHs05Ja1t40pgqYIS7pLamtCHkGqsI9hz7mccMaSKeG/FRMDmte7CALXqRwPeCutN1I
rzNKBTOy02C/WWVzrz5EetW6Dwk19YbEt62HNLZGx4CdH16fng1fsfXdFCSLr4+jf8FQabkf8pL0
nANPWCmCOavEDCjfnlKxKzRrZuwqxqhYtXyRsiRL0YfPRcRjIUNIxIIyZivSwFGEc0z8adGxNY5a
LuhDqp/GeKA8uSfVxbx9WpTv5hZBd+Tlwh2sMXXh8u6dnVObWOzgOzJ9PZ4tGRY67bcWjpD9+J1B
br6iF+RBu0X51D7G/7EAYAGkRzI9xgiVwozuLJ2aKgTArmDGkwfgV9s8A8gpiY4JM205F6FrYyY/
VGdadvyXgVS8k8H0zpeY2lVptaUmC3NDXY5RVfSvTsvMTYEvOED2mLMTMfRwgHwVMY23Cz9KvcBJ
S8VWIvfCw5ppVsTFUBhR7HlN9DCMkZU3B6dum6lW/m+wypFLNY8+fiPFnkiTBnouar6OGiLCg2hc
mmri5Chvg6I00T/e0EWG0eLzb0cNe9nlwJFPinCcOfu86hbHCTxUk+VZisvZ4NOjnaqnHRWqy+e0
J6OWf4S5QgOD9PkRFNDfhB2gcDJnhUJ7ImNI8p9Ede7Upva7nsooFZJf+Uu3cv7gZ3HRTlgxQoY2
Iwrd+hRyg6cPXWRY5eV8soQs2ntTBO/dtO9rMRThaXxHSPX3SSu2bd4xpvq/2pZQnvTtJJ7BprAC
kjFF32agp9b9/ZNUBwFV61FAqumcR/HpOiXcpJHMiDJWq8EDFiWduT7A2o8ChHejMscXlkkKNI64
fDxm31d/o6Vmk4bnzRrFVQiY80MgMP4cMjZIAUq+u4LHWDzlWillp7B6xp1t1eLS+8a1sNyCQ9EO
GwmD81tqJymoBylTqHvTYOronvuZI9GpNfPt9DiRGwsu8XHhdmuUJCUIHsWsL9cSDmUiowt80VvI
GnY2TAlqYuUBK1H4FzaLKDpXqIenh0B0/5z7n/Y7kylQIBDwP2DpUWriehu/WUvqomkNUynydgQn
grqqalV0NBHbc0/5E1BUWrZ1mHoVR7ohhs6+DJMiA3NcyBwcS80yE+hw9OFqGUpZ+GuVPjAji+0y
BHzQVVZo6ICG6GiNd58DXRoskqsFFHz0wR0ZiEuxy3jB6k4QAWkdsk7MpGFffP04pWWixnQxtNC2
Zj7dJ3/IQMAz7tRLbP2K5rnA6IHiUsMgWegCqikcVakiBnnxP540VzYIgqs1tFnrBlhfNCUyYEkx
x7AbzgcNgmQ291QKQNuN1O4qtCyAhcCiOP7S7GfYJm3sjchS9ZwwOlPy1w7mEVpJgx62u+K9gkIL
BERxI9BQ4AeH/W0AZ8wry0cPGff07R7tDceohEqsinikI1MEBKRspm3zMS9220Rm1oWukfLQqU8l
X71EaNxzGUgyMJkzaggVBC/utGDGfhv/0nLWb5oNPqhRZwXsH7NT7ggQvRtKBZxQZoJ1cHzA/K6n
FCTYxz8WR1Y1qdVeFgWiek8GgdXg21g0RKXvj/GtLvfNxKtre4nwgsXEABebO6swnHMu2X+1jTMh
AKDTMT+IheIrPoKAP+/J5f8tlPAPaUNaJO/OnAO0zUdULpGboN+ZhFVd3ezIdgy/EbABUa3FttGC
UEDvWGIwa7oHif6dSys5OY/mrh4iU6J0zn6L2a3F3+n8PkYQRLvUppqacH5dqAVEKIVzIFvprhak
l60REZknqAjLIKhu4UvDYrrqEL+Le6HgN89gyjj7DOvHL07bFFHcfWPJug9Q71JF4GhhE82z5E+I
lcM2SaHvr9mpo996jxDK2P8Q86dl2nSyTbFLhmRxiKliK4xVdUHbGt6rnaiYz55s1gCV9RmcSksn
ca4dA0TdiYse0u9fRlyS1FVNIgk25sBYR8RKs4pjlnRoqOJw8MSLLBW2YvWRzN23ardJUZq7sYlw
dlQDGkiaqIHipAn4aC3ZfCFAU3qjLu0vNgEnDZGNeMasNA3tpNzrcfQg8s8YiuSimw9lSDxA9MH+
acLaB6EB52abXewhcP1qq+kra25SfqDEIi9BqW8tjNFK2NQUeAhSZ4sKCXuO9AXgxpLJYZAqq8VQ
3GtH0Q2VYfWhPLiafEWON4UBIJpPKCQbwzIozjvNWALmxrY6d29MYtmwoWLDz/y9DOZrPYsZyxrL
UUwiGAAQzD+KeEZN26sWP2J8LuMdI43L/sEc1X0/mRP2ILrSdHuYc8vbnpVvp5rAiu+vQtJlV621
Lm3mOV504kVGSRB82QEUviqC43xFLWw+w4YK+POinK/IIJFBBEtkjorUgFjcslu+sz+sKkOjmByp
GQMW4VqMze1DTF2+EG+i0Ir5QA+FD2e5AedeCfje6elypIcCKh6RSGMXqpN9lfKTtPt//IHtGKuf
04xG0cjTfN25nibLZJvznm9+XLNGVQsSc40Ui5WM6fLFKOtrZwkM+IrZBkznZWmiUx36nVMA2O3B
QYfdkUuHQLsUikkTO6nzaJ0id2I4fvY8p1f70DYN4dInDDF4F8R2gddCl/Hf0GECvmnRCjuZ+33b
tq81jKU+rUF7bNG6l0kD0vP/HXOE23cm4pUyUKodbZRgmZSujX1TnGDLSIrMZ3Deobo4nWXxfQK5
pRypwMN7LcAA6sLAOTq8hv3s6Pl93vLyFI/Zijcrjlv/cICw+U2UiknQemYp2a3Fb4PLfVQHspoh
8z/Jgd4ovVJBMQuuENsGvSHh1mW33aSj4zcAa45GOtul6Vrb4WgWYiWVZ0FyNOSlwLQ+YKc/xQr0
kVNOs5yh1NEbhlVrh9/CaTwJcGrIDhOeyzridN+WSUKbdpmItA7MiTOPcOqEbgtET0gj5nSdV31y
NJmYvcMqTJVH5kDz6cRfGxRHwELSoO7bOoy4D86ota+wz4KHR3KxnU80b3mbeDbOnTFPOHaHlpbV
QtcNMjPFLotsImYa6O+91BWsdN3XZAjfv6d1jVIlBYqlW3GuLZhMMPKmuQtep4l0dLFym0u0dKlm
9oMU/SVCBqtcfGd/3Rl/1x/vF48wZT59GnRHK38yO7it1VZbFALXt6PABRduG4m1/vicA5hlhmuT
IIR1/rB1wQkbP0m8no9U9yv2GCGhuah4A/F1WZ/tB6QDXLNiiJ4YXuBqgv+HFMx6F3HYLPxFapiS
hhyjXS+GKok6NUGiJanMRIW/aHc2d1nSeOv/ZvXnP47GtS6l9tGtxZu4rOdK+rlprgkfGi/r6yW0
biNiI/FytXFcbTkIJN34/qhHPQ2UxcKFB8ZPQ+CIa92xSzVVATHzgDaAWlIPH2IPVLPMGpRVUTvr
V4fCwIUtZQba6/rbx7y5PV6FzXllBXwM8lY6iAYuczJ+OhSnxnt+J4ei7GGGahbegERqkPaeWUHU
0W7q4RmS25d8KJQy74CNp+cuJZBbRKuSh8SbTtVKM7Db5cdoXwrPsYAwW1mcggCd1oN2BVUXGqA1
yFVJqK2ZacejZiIGpNz57OqTIcxZ1Z80SK/ubx9dnqjxNHSy+DLcTS66erR15qYVbFaDb7NbLhUL
NFVbt+zvs944t4MUJ74Rnx2eAtH1bFIymBq8H2qAIylwdHjZ3qYMtLz96gLoKODjxYFT3VjwKJE4
hB34LEiJ9wBZJCTX92QeEzp2rSNTyJGg8KVi67tQ18947u8GJnhCQY486/JlJVXCE3kqEeNaDdUh
H/5Zos83lBNOJTzWwyGxv/lM5zqFAU0ifpHSqNriUHpUnOOUNh3bm8/IRsbsjp+6uUEifqE/OpIK
0gVCSwDXBAb0hYHKVGz4Ed5woeJ2U0HyTfrbjR3RSNnaVAe1nP9khVlpiby+jjPsXlq8CdTcnnve
bNX9uze4TxqhZiHZx/XwyYKh3gR9Ks1dFrDLK6Ad+UxQdQjI/CKGovNbn+M3ubbYJmrzAdQ0SYgG
xxaqfetK2XSYWk87MLvnQpxZlixWVrIHUSZjPsfdD93LwWOY8uq6iHKdjtv1ClXWTTSVlEUtOgb6
R0Ij+VEf7ZQwUnHDaoMMvI2yTQV8moPM1atmRk1+Po8hPU3GOMv3Rhe9cMUY9GRP7+2t0TvIptSi
sywkMU7p/jV8QYt/sF2o/fHx1y2g4D0xNESow35vVryHF4KaWOEy9u+Wgq6ilT8gGtbCFNy3uxKY
MjWKG1yzzos99vAdRYUM8hRbo+/L+yDi0GIqXAixCaPKu94HvrsNP5NVLy4W+n81D8bR7vbXoTyj
MFJmNo7u1LkPJZaD6c/nruJC83Y9CKmGVFj+uTKbMJO5AU1PuvB04JsuAmUWdgJVO3fxKZo9WmmI
0f/0/i9oKTQ1+Hl7JOyUSMXEvCfJTk4nhQvLhZc9r2ZLq2B43fw8SbKoQzy/XSKbUr6ViHkrF0Za
pbdRvHVgeByW8L8W8ZDoJ2yvQlHGl1cN9T3gGetX1USG9umZs8khLIidWq6uz1sSCxw5NfEA+LIo
6AbH1dTzGJLZc1/sOLmw++l8CWs/bFhB3bECnlnk7YpUF0Ej6lmhZF2N91Oztjt5pLi32Eqge5E9
3lF14uTCLWTd6CYXQRbx++rrg1ptXdQqpWNFpIaZ0Uf6U2JiLuUJgDo7tNrhTwl6hkm0ge363Zwl
Fvj+uXDNiYpcAvnsgAKpe08wlah3+jpeIg/sII1JPYnI6dKQsDYBIM+frFwKGgz6HDb+xX8a51Xi
Y7BznHma7XFE9k2WkbogqDKROu37O3STIA9x6qovnkKneDs1i8nvsZ8dg8zWQiZ31o5a91J9iClp
W22bxXayN9FBpYLM6JqW+KWDIgDNYOtf4zaUjGIsE0QDc7LZUiiAEhRUlECQQimGK9dOXn82tBKk
y6CZsccOtkZxL/xP6gfoe2LtljQ9MXVfmrQjvhQ0/ZUV9A3v0HUBqJvfspTi6XmgR2ZA3QSi/U+G
0ZkqHBXTGukRisOm/mV4RIsYww7b74UKnsNchK7MWAFckqN30wU9J3Lk+6GM34TQVCfa94xIS5eX
pNVnhe8e9mmjTC1YoiIiCOG31h7MZsGfvZ3X47dT1SvS2Tc5/2+Ec++QapSLOrdFaiedqV8yzLug
m5m8xgnB4x3O+Kh7ryjN7BccgJnTzWyE4FqJHHLmy8SGpZnQdskMmNzzf1jUFt1PUJ6AKt/vxeq7
Xcbws0oNL1qN31bfzxUXzOrhnQwLZCE2FGl7F/76dN4FcNc8pnLX4+OtQYSsebnAdwDhIbdUCVBK
msSgnAO1eRTAmUBUSHWGQ4qeqDqh6f7/q4QXP7vc06uW2Q4NS0xZU3C1avMDh/up06qiG+BFswN0
AVjIWSbUiIbJoQ+ZhFiH4qGxd2ZnPO8jzm6sRj22QkILfpJNT8mW5ZPx8SaetUm1XiZDwKaAwaAd
4z6SoeUFFotIYAnXald1SpCLFRfIw0xeyCjviDn0bGwi1gkXub5j/il77H6tvZVz/SXGFFGpeuMy
ZsHSUzqDMm/DXpCIHhYygEBIFQ+RJz9QgR5qRlIVxG70FBJ/3+bnhDMhedFhu0wasGxOji3sPvOE
hHjcvv7//tI0ih3kaIcStHzyiwDOBM8AKP05MQYmZIxLw1hYDBdsIvy1C50cFTH9Jb3yseyzKEfq
hjDHnT5wbCqCCkMzXjc5XafiouUy/uzSGdq6ssyfIEhE4KRMJCG7NmPQxsOqG/N9M0+LlBvxLXo8
nv/DHU/t3UsZpldYi6XrOmZmxt5QjFrdkY8b7a0RjsuHjctVqjhinIS3TrsV7NPsmTmTA4NV89bM
NPiztycf9seP6BIFqf5wLC2fZs6Fs79V+q5fZJOPHMWUa3oFRbqXrnOhWjR7FPs+dJlw7BQFsuC2
ONBq+oznz/NMAfbnGBUSbA72GCgAJ0UuNYTmTENdgzmAj+3S3Kd6mne1wjqEsbR+yWAF63UpgDYA
l/gin8uVv7vGY4HmptB/7c30sqaOq0WEgjBh3asVCQngC7xv/0ibe5ubLQrrpzKU2cWN3DIfq4tl
TknDgPtIciJfxdH4KGhgerZTo2Dif7i155C7gAe60vkIprGnwRvUZ2J+sAkAyZ8gkFJaENQ/0Chk
vY9hLx5LHGiqBNz9dwCgv9dD81Tqsl3Dth4VtaNmo52NvGtMTjw2f8Fq96AE0p06YyGMrMljhffh
TW9TSuKMXyguyzBMqSPl+Gd1NUNoiv9WENfJ2JuDdprbBPmf32CPzPeX3yj7eN3nF4qqvo8fPYz8
x/T/f3K2qEVJzrAtdr381doM1Q9ZHcR/HQoOtU7JCYiS+sg/GP2sT932tWUiTheJOTXJ1o1QNapz
++9/QjCwwST1a4NsDLWlQWnTUyuhkb4o516UN3gt+eq7irrHJKv8LB32fXqRCasChZR36LlvBugm
VPuLoX8BI1Q6XukwzKtxmyvnlDC8UjWGBvrpKVib0E03MbE/DvRO4Ex1c+q3d/wWHw27se+RGpo4
IqUU232AZFOtC+FfmTaNW0yVBX1g5+BxEZe5kfxBSL3vJDvzreBWQy9wWN0Er5va3hBvWRlPFkBL
k5unYmy3u/WbWJ7B+I/Ee0RVV+AbxzGCF/s9BS8Xs8LT2xMNFB1vUojIDpSLatVKwfH68TBwfcUK
z4GmSqR1LdRLFLR66M8F1BTY5g/8hRdF8Vz/0At+YQD/WUAcG4vkKV+ryU0YVbP15fi4i004MXUc
50kVSiIClmf4z4//FcqCPAwTlTlcyMxc3x0Dses7Jt/4hFtT/ErW5c1q0VbsRexg5nItP2hnw3c+
3unwYvDfum9PATAfzuB97wKCdSciCTOMuGAZLUlo0wpRZl29W1UgZJLPXs4vcKpZzif9M0jOX8cg
1b7w1MRHxY+kwG1evhUBIj41KMdS3uGvsKBNkj3gw02gLRxBRmPTWB4tUYf2f6vMvj0N0frHv5C2
RAkmmzyH6Ws7KUXX2VATO9uhbVakDYjNm6m7Yydb00J4zf1/s5IxOP/ElqBCS9CQtEK5iA1N/v8a
RoYRuAscFueyH0CC6I9YubY5iwVmcMsRyjWqRsTBFIoytSLZsRW8dBC0Ok5tjTPatx+eSIs41c1Q
aTQ/vKknsr6Xhpnc186yBqS25JuL8q9Sxb0DeS7fRrfh3+HQJs5ykjx1mlo2PsSq+JN81OcKXLK7
tuncY6yi82dBObSi7dBZFdXEllv5jLWvbwINproD75LDDgfJ1HimHEK0vmXEZNOvxxWoiuvcBBq4
1AZPrDef94GzIKKu9h9pMP3BEiyS3eKznFbFPcrOFgX9zIi9IyXYJB0XS8bFs08xNzZ6jpN6i0vs
9OzDDZfTEFd1x/pILvQGKK68+/TsdgbmU7kCWow/Di0/EB2zBsFPD/+ZY7DtNxFyj9lzCh/VC37B
7YTSJp71IrmQTcUUyLh5XM1fpeOAJIDnYM3n3tuaqXqSazYii1VYT1R0CxKsmdTBI6ZtfT//JqHt
Pwnd5mBX+hfxK+TioNQtlO/Tn04eIW9s2esAM/2rLP7KAs46Abg7a0uT90HyrJC7d4NpWqQINBUw
wldSjpKrNPhGS08vQdS23kafh9sg39B5dJoa7M1eXeArkq7c4r8oWaMubyIEPu2cdnUSDOqo3Vl3
hrSb3gh3j96IQ0RWr0juurbAXLrDk0CYRqRpDGRGdD3dp6Eys0A6VVzqlaExhyli+IHHeE8vDRLA
0frk4ePod9U+pVeAbDZhvHBbb/7dt3xJ2jFoOXdmZ6nhJYs3Sx055YLQUs0PK5xwWsXczFgIGOGt
3HFfUqfpap1mMqx/b3Mi6FQB2jIRFpybySnEElC3tQPf2w5VV9XhxoYQiav74qFaJTIhWtg6tV7I
h+Zk/Y/SuJkTkJFg4FZztNtmX5ZqSiT5PmQjgbJE4gbOlOewZLrpwg3aaKeduHMjRolIJn/Y6T6P
DzrzATiVokEicOEmv5u/1TGrkr1m/UGDwxCYfi8pRFGOEV+a85r8gHfdjXMHcAfymTPza3xLmi/6
S9yMCU2LPTon/suRQcNXXXJ0v6cE6yjqvckkmtYGgLYZQb93oggdOktlTBzIDDKViyTqQW9X+xxl
i+UyTohRnaTwvaJlLNwd+REaRnpcFCpe0ewfQvzjMSYfY8bmFpROfzrEYt0oEXReBO8WQwQctoa4
/CBL3J7jPQO1XuHPaRzye2WBzKyH+adxNjfd8NlgbBZDlZZbaXrgcnDuIIrGgiGLSf5OojH9ypJb
RXze8cpcV61lXyOx316I8XqlT5dzXREZqHAiVwc5HZu3vTIFuCiscj55GHLc7YWIPqAgt0lCJtmi
ieg2s3UCogG88Ug8sSwZpHA17Vaah3RDtzhxG2vhm13wdTgtiIWQ3t0kId+QbW6vfP0tvY3jGZMd
2CkkX36mh0Sl5u94FfzboQNPunqRdXV7l4LeKXg+XpOcUvhErcEaml21Z4LyRUWzKDn8IN8cGJYR
q0j+RF6ESzOIYxVvOdo85A/rT0VwrhfBPUBRWNV/l+/mPTWg3dcrAa1YtJBv35xa14rx/420GSaN
HTIV26HTgD62EfwaxP9sXMMtQ2a39O6k44lO1DQQbB+ZkafZfTi08dsv1hW0n6CLJpT++L7GvQ0q
PL/BKy4i+sxVC9aBT3g9vbjcz/KRlo0FDH+51U5BmUrnvHyTnZcPvIAvuzvOP9gfRhzuaCwdidSh
OCT70TxGXE6FKxNj5LnDZd18ioWgNiLAX+k2cEcolMB+iD9bTIlF19UgFghaAHN2VetqFDL7HIVp
SBDg6TyGxTcB07agtZTgy0eRbPCg01qAmodOAeWCj9DP5Isl0aPGSc9ljrbXTL1ULm3oh9QqpHoI
rQHG1OieqkDcz9x/YNI2atVOKeduSgPVWRkOVIEsUrBkWdu2j8VUnN1c7eBapHSaZf1imJGJuySw
ZUhbPq98KtVoN31f7iRxQ/AEUACk7j5QTBytBlsKo0gHMPPw/L+GKy7ZTMrOL16FRrdeY0SVCR53
qivz/H93KPc1THaFuYSBXjEJE0S8IMFQTH858IwP1GPgwpZBFk1wcPy1RYvRyEQ8TjcwDuplhQHd
3Nc5dF3/LUtrC8BxG05VxiiS1EPN02bDkMnKR2CEln4iiQ+wlG3yrZQ1cVYM34Wp4WisiCd3GMfX
l/qnZg8+08v5t6RH+15pqU7D0ZaxKJxGuwWl8zdE2z41ufCYW9Fz1SssSKEXCHCpcx8oJk5dOnVo
UUClcuzeBZ+qi+PD+s//Q09n73D1pPM7l2f8fVrk4BeMgzMEUbBthaUDh14hqqMhA9bxtgSd7njA
I/NdxYjSm/CMkTSMxrG7LoL0Gp2orbWQAUfHydb8BzJnF6EBLMBwL1ZL+h3tMl7teqoewvMrSSsI
UakyF1xZr4D4Wgv4lJ6Sf4gpkxYBUZNakd9nIW3r7OVDKTP9l5w+GSU66ObhLA2ggSofJTFywiYY
jMYm+F5ga1ZwyLLkbqp5YkJCxKmlrI/cwS0dSWuPWZx6FeOaGJiTHV+zPvmyEGxAlAQA/UzaNfyC
+CU7ISsz9xqKBY8sc160h87AAQ00Bb86oBcdoLuncQGIBbCOZFANsMKqnsDB8rNqNJL0UrjVrWag
tnIu0elaRPzfCAktxB6SkPbq3ky5bFxJRxT2hxBiyi4yVQ4ecrXvfesdwE2fp/vqUVn1LjjnoDS2
xa2+/s35b/0fTxP3tjudyd+0YLFsi7elGHebKpJEjf4cDjDWd5eL0vXzrBHpif1auMnqqrU2Srny
gy/GLbraPjm7dtbnq9YNMMhJbbCMUz0SJuqQj87801ARjlxk/e+JFdYsTymLMdQADpFhlJtHfBQv
jOvnnPYIApwQrVvQHFqTSL+LKAx7qsrQviRid5eqqoV+s2cXgMQRzdDrW3pbiQ2rU68wuJwwodpq
S0g3Id68WcIMyU4Ck0MbzxTeS4FfFgLTi6sfjX6UQOMoUyuKWiPsSVQelNzb4hm/epXRzI2t54ag
JNPqPmazuuNoRwdGj3nMv5qMyzVBDWqviBdPvdlGMxcyaxzdHt4bBwYaPgK2goZUVpkrH98DCLvG
cdA5atBiAjUFmn5uFh1WIQp6h6xLkXKIaeM/dUup1aY2QU7TzwWBfYiExB3inmfDBRmbfIKdxFmt
StVPVWYwX1Elz0bnPlfwQPv3ngRAkIRt42gFBNw+Q12rlabkREhZVQyGWW4Lvm81KcTl3DibEn91
A624M+2fsUPHU6vOe8V/gTyfXTPq2Qalx/Yz7XdoxHNsfv5eMo6aYFzPAtGpCLApXhHYMu8YTJ1O
d0dUhAdH8j+bJ/CRlSz4/LF3Z/UqmZlammD0Kz5plNunsTSXjQOilIpqL51os3szbvdUQLIsL3cv
gpTIdKaTuxNJyczORll+Jxx4YNZIQY3EwI27cxPBdeE2ia9HP7aLDMTaqlNfVshEGUyRcg0C0BJC
0sWbnPBkpjrZQxVN0diU5jKkZ1xPlWEqN98UvcZdETLuqfnFq/PyfwD8wNygEtJTFpjv6Ml06dC1
/cPW3ha+E7HDFGbydewf+vquoF3b03i3AXDF9jJtQuG0Y8H5iwoL2rJdbTh4LLYLWWPEyHkfGwZr
gt4QfRvl00FpVzPw8ZD5GmTUDyAUbfA2tsgexe+Vz0PAczftGYAOFZxJKFQDKIdweJQSUyrP7pGm
Fqjlid1g2I5rGROcPTzVC/BSQewAE2N/xs4WNZK/L8Kttfw3WbBwbiP47anKF+ChH4MG+AHdrpCV
/rYEi0MMeYnP78ksh3WhwVfCRArRNSC0lYfTS+aIJC4dk/x4Qv/m+fbjh5sFAmY7jvn2EuoD6qWt
H6rF0WQ2ijVQKg1AN4xuQBF+51e3fXTf8Jx+rPIn8GPVt3bzdqF5zt4dR1oNb2P9B47l5/EZ7Zn5
q9W51DEme979edoFD8CJQt9H7K2y2PpAtxneDeyjQqFsf0tntYob/jFPQN4YYrshx5YMTUSuiBUq
8HRtOF/zjJurBLJHbIzIy5fZk7eJvN1UfDkacawPQhuwafsEjJ9GhQUk01dp7AaaPLF81Mjkp1CK
1DqMFYCY9mwyhrOVmK9wqNwZYgzxjGmS4kXs4EAfUPSeIc0L7+8RmxrcA8cqDlltfUOINKeAIq7/
Qcmwa5izjvVL+Go9Qtwa0tZPpstOkBM28BKY0KNB82ZSqTYv2+pf3zwxbnItfeAPGHdBdYI5h5IY
7I1A//YkXGsPlhmT8Av2qshhjsGlec7Go68e/h04DmnLZkA7xzpj1tzqH2XgAXPkMZkMh3jit/7l
1oB05ND5XBAa0TZ/x1UfeENRrJeDXBXOXdsfycGL6TlT/CGyBO9Xqksd+diX0F3fI7DWjxu5KLmn
SrKhMuYyL2QjLs/ZlWNUB9lV+DByRamE+vtSLrL6XTVRI9hbC5/L6fAvCzAVtSD6jukJwRl04eZO
6CZrsyUtbIv3OyMlbIoAbfBqgAHukoutRHxOMnrDldCpkVPFNbj8bY1B8vc6+Z/cDiMqV7BXIeCl
ooiNdke91xlavyJUdjiqkDgL9NfzqGx97HT9o9boVBhHp3tfXqPDWxh++UUVtMr4yI2Vz4Yb9dKp
5k2z3VBhHNBla9xNXd6inc+IE7n+hGbZvnnVuVMg84UxoVDvWnXRvnVWMGmXGkDsHRIpI6ce+jqO
0UlMEAn5/NAFfp7VFNa3gqESF6tQM0KNudxtQHre7JPzcA6pDqjIDZROliJYTxXqr7feM+HyZlyE
D6nz+kQRU3Bg/u9mGBGNQNEYn3AizOKrfTv7nJUKpAQ3b9XHkfyXyjbN4nCwcVdV9rvKj/xlnFEP
VkYyGCbYMrrHvqmEZfGmoj+4jjWomz3b9uFUb9dk8KytvvH+n+iIM1nyuZVDdmOhP1lhB2ZcBghZ
8FWEV5nFHVWShezNTwBS6fskvkhazunrZ56He9xqzkzDqKmyXJI/NIX2P7CVdf+HSbFtNm62q9D7
PZSPf/SZLYha2ScsREJyTrtlbpvtTTvD0RZqFzhgdusQteeG6T+736g3jjSnegEil3QOmrXthEuI
M+Bn4qsQqFRovJK0Z7Ey5xef/serxDnjCrt+1i9AXl0KusR5nWaHxLqJFp+8WXjeXdd9SeHwdONu
YWSb1I58ioXP9s0L/LdeOqcz8pWKCKs+Tb+Px6bs7EUQEEqjkTTX6tlkh5nBkb5cjY/1PS8WSEza
YPJfzp1WCmZQatJXC4HAYVN5OMMJ7lAjue8671otZOBc4ADo/bXh8ZzDU/4srF3EKdNp5No+9k1j
d/f/5MofgxmM19WdLhXhat0qm9gFNL5Po890h0Qg/Yv9ue1J2v6K/8cpv0KqmAMbZeFM8eI+FWR5
3D/aymQRyIfFMQ9MqEPsepJzrs3Q6Ve9oNw0aHwSfUuR6fuM46NA45ayNPLQm8F2fsl1Vs8QauhA
EWQENEgB8K1gYB9RIZhMdp9r6JHIw1QBfufCaGWw0Jjq1FFHe2hBWKeYbhdgaqqQA/1NPPVtf8JR
RcqFuIIOu3Tbzuy5KrB8NWeviSnOEYXnGXQuIKC168lqn+5cW5VTuYsaZuO5k0Zyp9Zs3LTvacP/
W8FZKYGHX4iCcT4FRP+A/tE+8k9QOZl12XJSGC4OKYDO9NUKRuUaks0QFJrtspoF1IXypZx8FJTE
039EG7QZaG425xBoGteq7RGs0JL2kmGw7orLR3z+3dPnvamndqqw341qIavTl8IhhG5IzFJDGJZn
88v6D7q3pFcLP24x+s0ka5keGVhuuxZgk8qaNhAPMufKdJcD/23atJ++UxefpnKuaWzu0LTqgeUQ
fxjb2doG3+HOUNAUKla+CurmBHRbNcvPZ4h/5yhYteOiMR4vZcWBk+YLI9tbKPhnlh/6F+fuFoHT
pplZx+6WmturdRfLndLwn1VlNtMXkS/YgL1Lb0AF7ENPYRKGvmv/nexOnZ1tzFxytSv7Uhsq0Jlb
elXKJhkb5durIkeQFY8wpc1mfOXUlkK2ckeVnafwvXjZkVXUDW97zRbPVz5j8Hf1fxtwZn+QpQ5g
XGlBMWz7hnRbYpL+pd3dnTH5eZDZq2Idl6Zr/B0fxJBLRt2JDYhF7zPImcw90vvm0Kijl+BuxVXy
GCX4h1ZO3emo1VQULXwdeYRpPeuq20ZukHx7f/GeS8k4IJ6aMVZQCNSjy5uTi2IRF7pqdvcKM6LA
1rSgW4Bnzwfydq6vC5E+UItV3vqw2LfMEDscuhpBJweRa68feayKI3G+dujpv0ktgR4jyxEsUVe9
KODLK+sZ7DHOs5WVZcGaUeV/pH22WjJUC9FdwWY5tyWLYFvRsmW0EFoUgxtQlkOOVZmTtlbX/8IK
jn0XDmt6fhsgzqDQ/NDnoaHvJdFYyD7L+bkNoGUmHEgp9Vdf2H9L77psS3Ogzumm0EHfqkayPl02
AgsNl63MNFtMn3YaVUBf/LLana8rAY9UuoaW5fvokstiNUSZLsiZmG3weXo8e85s3oHLfrU90zJy
NkyumoMh/MYHoItaV1HPFTDqJu0qv6cwldD7szoNts6AMoYAW8ZCClvxxhz1g3zt+QwQmIMb6zH9
OgblEwYsskcsZ8V40C1kyOO+aJBCDVa++IHk1kAirLHoL5sI/aflso6VQXNNlBQPZGIiRI0Pnu7m
N+ibQtuXvddphpMYdwnBsN9q8KEt/ilLPOG70NQLL1lQ6GUm5jQam+9G8FIqMZi/48yXIOMlyLwy
GvPi58FQqeRo/arS1Ub/LUV/AlpMZZcTmUYx/s88Ps4mGBOwL4jm8BtV0BdvNbD9322GX+0Iwl9V
SZ4RvUON3KZ4j3VMR1grNsSRIEpLPqL0Goddr2gp4n6c6DbWJbpMfpxMRSebphDDdQcx6h/oMoXb
/htJj0lZ0IhEd0/JTDeqSTUTAwTucGhztPvHj1IGmCb6kyX4Lih19gU+xTVCOB600tHLwH+ym0cs
pA6AaBVgy9y0JlUHBA2owKDB0VVMvCMTdHaOcWXT66if0Pt+eEbTb/L2QP0QwdY1U09c9oIwp7PO
Kmpl3JRQvgjIxkt/jpS3ONcQfm9qxvqZkgdPtr/qVjT7t2bn6VdPgwPAD8JNeG3afGvaoNzgPOas
OTbphuwtmckwB+BjUufIRRz1nJMWRMIc30lnctXc9tkIPJJnXM3PHblu5RBJRFTNaNqxHJYkC7n1
/a4ecBC7x9ZVSV6BHU9DmJFoJ1uKxcGBGOBncnIvQh/KD39drTINr2VQDDbBzjSZJeGAo4SUQ5Kd
SfnLg/ILTiq4u7oj7aKhDVOz1ft2OWrT7Y1ll71tAcBBaNjvcsnDzc7nWc4ABQkHD+G5gn/PNTZm
domut29aGZSNMWVWT/sEURgotyem5EsKwLAo09nzGFF14t1OGufTqn8Y1fH7DSqmhQhJ1bp1KGT7
JpFixoEVVIOP8vdZ6PIyShkdfvKjJjzAcUysSgcLvxV7dUPYJe6cqlZ7AFYcDN4JqSfb/4PWVNGs
N9nv6+eU0XFx91b8FJ0xFogvWdR6ZKmg3vWCkgM6RpNkcq/Uj7luuoK717z/o3YtSNa39OxwLzzU
8lh/KQduBN94jVoZTwWUa6I9ii2+ayBKAMCs0v5MWhVBa3DlRPwAYO/dU0reR1VXjJUx0/aofSsN
fDlay6qyaklAF7lO26haFXwkBUe9JSz72iV8C3tNIdnxZAJai79/x/THH0nk2n6P6jdP5fpoGHib
A+wxhNTZIOR7eLn3Gf563ndt8d3Xpl50kdfBrzSOvvs9UrVxayNv1ZjL03fTXW7cWmB1XUho0hMT
1c0YL1y4sBM147J1sbl/sbIrsMJRKRsaSQfib5Osc9nvciM4XkjwQloXm/VMhifqDt9v2e9Gpxfu
oI5ioYvgH+5oZFf08jusDsXpKjHMahgSdMrLr2TZJJhm9Ez9wPypcJPA8A0RrV+Z4yCtEHk7EH4Q
73g37DqDmlN8aPxNh/eAVbfb7e+mwdaT8AvTIv2qV6eauIFFPC2eGs2X2piKaSL7OywWMxNZ+BUl
dqnbhQQ/tjzsvjFHmpaKJ2cVBuvDLx/h/9mEkv+FRE3KZsq/algujT5atvvxuIFKt0W19u+zFGua
X4hO+asqGYTDn+2iPhI9LVhg3Z47CyPkI3wXqTkOM1DS9iVd1rIZSzhHblObv5AWy/sbifMZYvTq
gtE4C6PDLwPujKJojT7FtfCRyGJ4AXdLiroBEwvUj3MJYH1PdAhfq4sBixLqlblcmCjKe7exMtrh
Yd9nMxVjz51NYXlE5gBVuBl36+B8+okJC2sTFSTW7UDDHpI2t9/xDezEn45kiDyUM7dOvdoycTmi
vR2zfU/z0zFQr8bmkV22iOMfb/eOfv5suUmBJQUClvczMHipm/q2MAbaqrBHcAWUTaAJcB/KjB31
MNLCzx03qqqbBfDLS7bgPOCfJb4mb9XAzfjhChO5OOr/ZUdZFohBaXhzuNad+6EVjDD+lJNTP3ke
N+EkCSQag0JRqEGKs/sx6RE33WhRGq+lKmK/juhFrgiIBmyGi+z8eIvgxCjqIxUtMaOl5sfE/9WJ
MmKcvpDXrDkw/hyCKwGNz1rlza8EUZqbQntrEXAIZ49r5DJ7gbVXXU23xJ1cmUblF2KuRVH6nszX
hFJDSMsHy74K14cTZWcoFwwjddgzmlfRGWakEftNqgBZrgbNq/rsdtwFS9ypSVB//mrF528MX76O
MjOtRcErB+qWc8UC3tsm9ULTepPbAil/jTdIvAazCkGhb2v97Db41FDwk948cx6S7dA5RMNCc6Ey
wX7qTetPglQxY2A7CuAo3eR2EWznQ/cZjjxyYH0P2bwQ5VHOm9pCyVyaRXqA1LJJxLpdLDWTD8Oj
4v6RhrpS+aaCOF9LRixP+uSXHKzw4CNnY1OKSZtV9JT9Q3SZz1LDt4GiMQ9CMGdAuyygcugZ3uuO
W7p2bBGrUp0BpmydHdy2Hul3mL+X1HJLyE+rDjgNad32OrGh1DNqLWbp2GCdondo4fdvHMc6dwzY
sDiq8HNkJj1+YP20NMYaBjdWJ/BravWSEvrvzz2vufxWxHBt5CRHZ6j7R7I0/x73UwwvEj7lJM1g
px5H0odJl7+YYLuQZrZDr0sOiM2WBrJA+403vNUAgFZOozSyPAytqvJfp8DRsORLkBoCgaVxIrN/
b3q77tEarWIwhyaKz42JIpEfNUsZvFd++66pEFrlkSQpPO99KC+Q1tesCDTI0KZN+rdmn359XKyc
d6D3PiwaBiodXuCZxp5n3r3qChuajqeeXKcZKOyY08a9pE3Os5IFM+03AVYr97Dfzc0JF0Zh/eXV
O/SA2sbFqVM3xTy7mh+JOOCBZ8Onw1Ve4lm+BKdCmiUUgpt7Zc1M3BW1iyQwad6BwqCt+wmW4gMv
FKdumfbFqWIz86cSrixeRTXPZbbreC5VeaH0dNreNUH2A9CQjdErWC4Pcv8Ymhrnmt6zQgAkWGb/
L78r6U2HI2vLJkly9zJQc2ubV8UWoICVkxF7Ij55iGShQd8x4KlKNUeOehilBtApvw3yra41+JML
ZU5Wts2DQDZfTFmmpGg1ONk8X1Fv9172Hmt5Iyuwpu7hvs5UN0FPUsQPvG/yP6Y+Pw+datZSkK63
Fil20RIvHe5VvJnRCjrZ123hoI/08RC1/XQe4EDStUP7OGwiu85sscdZcAAQmB8DAnJU2WwAnWRt
u3/0XqyxrPc4Y0BJIEIoMUZvE4xCDxBO9qN/zTe2HyKd4ftISn1wAuGD684TRsNa5xv/jA1MTpoN
OjtNinq3S5q+W5eW74rtjv/7VAN7t+yJ7FVPwwK8sJOY64D6rfO4rXn5x2acSyd579jKEdUDx2B8
eKL/aCLXjmOGUigya0tXDIiHMtHfLjrsj/AO81W6uxroc8sy12RtKMBFRTR0FmdTc8Pn1gH8jwnG
7/hac7tUi9hX4a4rs0yqW03QswzgGrr9t4r+otsGlGhHBTeQNHDO1HO0CVx1s73bZnzIqbnI8dDc
J+a2b4OEriPIN74H0INk0u1zukbla4gG8eegKCAP7u7kG5CKPlSbtBX5aeO/BcuOlwmJAhpA4kkn
wHDBJ+W6Up/YxH8si9lhnqkxtcDxNKYx3/Ohlenv7VQrFewz8J9mZTc4cZ0U2invI/yxProgr8b9
a62mhULNi48c6QsNc2IOHibdJnrjRU5d29PKd3D0dClpq+nA7JWqcpYou+/kbo2buR10P6pgq7K1
L4jIH9J8OiyIcJgPXDAfvfKBipKZYb2LrV8MCCr8cVgU6HWopyD6wnmvUr6InpGgs+tKBKyH3xUh
lAIEnz8wPcWRIbeKEm9j+WtEglKWSPLMOHItOJkxlDOY5BleW2mry88nFV409EIcOzqntRIDJxFH
HE5MtafvxeDuUuZ5wGgkDXhQ9J65VhIxf8wtSjTUUuBCDFkCc2bGIxriVW5VEI88KuSjE424VtY2
+T0AYN3yHwzcWFKkBGxBrQRvLoeD3KWii9mebr+oGapBZTsAnMAES4SYwe/QSdsU7dmSOkau9KKg
IQVYKYTSORh/guRHBT6kEWGu/MrSuhS8ELgWLdf8m9S7M50ueQcz5MDunI1pOL4HhfzpKfmFVjtQ
ogMRS6P8OSmkcyQTSWPiiRqIOjK9Zqz1WbFxZREscj/B7YaSihou46o5d0GL9G7ikOqyAOLY84Q1
x5tMwxia6ajwVgFEG4eVqBsCexXX1vAisMU+oKwaJBYxwGP7VBemY1QfAWwQ+tXRCuX4eaQAiP2T
Xc8lAe/gbXQkPj15fGUehdZ5IZScAs9MlTSJyiX9e/hIwl4QJ0FXRjwIj5zxzHHNG+1pFFK3Wexe
KBm+8gQ+ErP6/9NAOQHZ1LjMJwYlP90pYo3HxWQL17d0LRY/8S2BaE30hpSTyQAOmfivSu6BjfHX
NMFlGffzorE7/MMDnkDDN1rh8OEC3AkGVT5g6BpL7a+BPExuU4flI+0n0s5lzX05SlOfCiSpjxzs
PBf8Pgup4YHjQaVRNWqLRS+TFKNBup0ae/3183MvkG5KWkM3mdycUuM2JiykwOUbr7rlv898mkWM
tsX6tdJ+i/aYWcejI2Kq2HIMESpPnwr9RO2mjZN7N6HbIIJHUK5YIx9SaoBiGcJtmuklMUHrmy9G
NRiEIg7BboNyqS4bt1rXRi5GWP8NsdTZaAp0MQ94v65BmxGWDPp9Yz7qPXuHdzrimBHaUjJlegcr
DaTPIXgabB2gZrLOfgdMSXksw4r3NuGn7rvWHenkvJnRxjy3UZg3icOyIz7GRxzkY1xzw8QTZYwd
kSMLyWHCiSp16hYoA7Up/x22ROB9MWnPpJDpgMnwQ+21NL7851YRFyR9pq8XUnlafvGUcL2+q+qU
HwbGoxtZWfZe8RUZnWOYrofB56lv4nrY65vW66bgVFR4DqiHFqEvEhhfcNpqS1fPE4OyG7nCeP+x
1Hk3bNpJsvBJ+jey77tSeTfYG1QeuEEt8oDyhtd/slqCy2YS8yFY3mCeRMyoYe7mwBJq/sPh2E/w
O9CpeCmaeAT+rcbNM+RquzyUq7zppgiVNtk1W43Tl6uaErbdlXC3nG4x6w+77hziAeqAYIL5/RWE
TKqREWizfVN2rzaq4Q0KUwa26/WFDYUwIa0e3YBX3Jnka69al7bEX/Q77K35Y4jP9TXhdZgjQ6TE
oqlEmy3sMhCN7ubPBAieb87Tm4S6Hw1cQzk+SYPrPQynpVGbBM0RGqJHtv/FKd7vx5lFQErPeLCp
Vqloi0hxtw1sdtb+6gr7mc6GKY8eqTVi0QhrKqMjPlhKalKFqZ8g6+r9GcLZIEjcFFaJpWUSSrOO
vbtsvHYfqb5Dw1NZvKsiSGiolwZubC3ANsV8B7WzF2vIsx7Gio++bRpsqj/BUAfsYPs6pcmG6qr4
swdvrPMG3ue5MfBz0hjfftTF7lQOvZPaqKERtANlvPDAFACtGxPRhqyNiJPYQ6e8SKQ4YmsbeflD
6bIcX1X9SOXXHQy3l0vaQyxO92eDjTzifRQgsJcjxxo+NZIxM8tv8tcYjKLWhjpebgdBdDCGSK+b
tt15fAL31a/RO8qyLzKnLzDGk++eCssPKgfzBkEK3dEjGHcnS2j4M5v2hznXcAWfr9HapmATBQe2
U700ue7zsAc7I6dxIQBzywi6o0QuXqMQO+XHSuRWVpZ3d6lV7lULMjjtWVXlE0zS1dPEOC51RQfo
j3QdG7uGNHP8QtnqWdsBkbapDKZuJpHu20M3FwMsKWwOzWgo5lhoIbdqxMp2a4Ve9vPxZgPEIkFI
JhWrL01m0VxIbzgrE2iYNx3wFLm1wxTtSIwJ2QCygDZbgWEJ0QAEnfX74oGx7Ddygw3Kw5a3Y04Y
SPx1yhhXlcTK8eo6hK7+1UuXXjkbZZSiisT1Z1g107rdy23lvbt6EOjWaHkpx/UhkBaN5ljWfqoM
kHqHHNxKPzmyEw6dGbm/V76X28ApmgrhWqTMGr+0tQ5zjxeBJIydnKKNdW+FVEd3jvgPGTBJtGsF
10eznuIGZ5HVAHIRFj2S1b7NrASxXVcIfTCv/3a+eBBOb30VXEsCtA4KgnkSHOyGy7WxqNWot7H8
fJlRfPqll7UHncYE051xDrdrc0to9IjUEc8fRy4unyO7v3orGQ3MsjxnsrZaydQNl07pyOFgm3ec
zLVta2BZ3mEvapq6EUOYnV3rnXO+WzArVATXVTAw8rr0ZvQr6j2+aMUZjUdohcoyRmWRtcI0GwXh
Oh2bKWRG1CbFnoDqFJprAPdmIDKpWHbl+1EhGrdq9zCWLA9JIBp7zrVbLMVme4N6Tf/fSG1lVze8
u1cDLXUXrQWsLFu7QlePhc/QteMQmsfDnZBTF27JuJ8NywR4szGNdp2TZXQH7hK5pJESuMknRaZw
1KuwbxTR3RWSJl2G6lRTmRl8Offs9EOCRTiEb3RSgU6WWoswQbHscVMIzICer8xt9IgtOTzpGJmr
/D/1wbV2wPk4oIn9D+3rFZJ3iCRCypEMbJj6obUOTDlFGpb3EziFf6CWU+1I7UvzQGYiRpptpKSQ
c4uiCqJiWebyc5HOOVFKXjcQj/5Rj2rRhl01PDGxBFHETSy1it0kR9LeKTuN6od3tCYZnD2/3MkD
deYEAKBhaIIc9mm9Xyc1IVPLgN6uIqlE/Cr0SWK2GU+fOPxZjBqluKyaOZZPBhbFKmU3a9fZvxD3
aOZpHbloMDMf7hpTwP8pMYmM7rsTr+QkhSwTUR9Hq0EJazX+E7mBo4kJfCJjRIa7Pa5osJaOrSzV
nywDYoSUy0tg3qNKHDdi3QR8qk2pbsFgwAAlCJCmnx7OpvDd1q17TkULN4MF2rfd9dLXJnqB/WCA
uqTiMyGXSsyXfD0/wS3HDexePvTYKn9Pb+A/BOLZVhfxdTb04aJRksKyVYQbbUYPKsL5Fvu97SMp
M66OERyXKYQJcLQOhLZ8RCJ+v3bAOyR59+IiKBl0Wa4jxzBX0GF+2bMF4LhnUTcUVrdHsswcVdmL
o/z7pRezKUXz3rv9Ps+W/XSYTdICqHUYP/gPPoXJguKAG97GZ/Y/fUabkBJmzQw58gaNA9j/k0Zx
33sOCjL9qCN40SEhJmca/bhZUzsPguxjZWiUHdnTFmCdC+XoXlGSWe3pWvjlkUYz1dPztI05sjAy
XUMEhoRi5+kJbrayg/PF9hdhiszK7v58SefKkgyt22cobkRhIdUZn0RG87B3fwGhaC9sJFp0/mRF
xrpBKNr8YMELm8ifwfq9pNPofZbMM2pD3XgnLvBnGysbDS6bviqupbJ8QGIH0st/Em+cYPJShmJS
rvT2at+bLENTgRfHVmfD23mdenUJ+OnH0vPsKAwjs0eQGh+nvIOtJOzjQd2SDmQwR6ukYjJWnVV1
sxNhBAl/FsFTW/LB6MseU6rxBvQVGKQOnKvmxBKoHK3kgBjsqM/NNdfVsngAnOt3V+YTiUQXkMsp
BsCPIuiq3/JIM+SqbBZglbAFrZWuCnzBPDUxnvGhI7w7Uy8eBlFQEDmCLTmoaMoACdfG9A0BiUCs
a9yg/fktLwOIc3f+39j02swRlVyn/fUiPw8IeRGtL6eWuu3v55sn/cQpE/voyyQA4p1wbKmS8qbD
PXCdWyKVhgwehNM8sVFcmQpr/3KdruND9hl8yfp17+tSxjgsJ1fSepSbHOwSLrdbMka8VC8UXV2C
Un5jqhFU6P5SKbEOkI3eRnwII4hVnGU8+0u4ygf7W4qtoHO04TtU2cDPXSNX416pyzSCdNnRdexa
KgBbQgN+WQpTGOfswSjb/EqT0lb4E33V45DIRNcq8l3jY6m+Z3qmZgWD8mTXy411scF3QnpJNLsc
RdenQoasBnMAa76iqwomu8EeaJQneGgA0/77LdKJUn872t/d/pYS5TZY/Pz58FoYx0FwCgCmBoLL
B9lqHg0KODbv1rx8Y5WFdD5XN6ubXb1aNmxGNdZs8+XzL3Ild8rmFMTaxheExvDwu5Q6j5bNJa+D
dedo7vNBlQ/9m+offCPVWQl6KwbM7yJVCDGRQuQGpqEs256xeWFHadhSC6WP8RdIbMy/rzCL3hSA
gbkthKgfiflO1lm5ffHsN1j0HMrOt0nj2zyE59Pr3tJhDMHqJ9neWmZTf9ASjvtHOSrzrhotIusN
QCuDBf4uNtEWsMu1eGlndVVHBFhWPSMfE0EEZSgj0/TZK5M4XgwhM01aIo6izpUOx8/eGiO89RWi
iBKEcUkS25OKeIz+eaAVEwGLqJFeWAiVtPSQ7mBEDDEYNwYAUSfl7Lo6DYzvjjnXJ2B2K3tnvyYt
94MQcX1LmnsjGs8f8Q86FlmgFtUsXGPHCeRWuw3SRXZv4pFCS1PlrfGqbVFTeeSRcyxeAhkpN16l
b+9JRHQr98bwH9OymhBaToSYl1ypHYZgYeRwmNEjAfFHTpI2ebjo3WUy8+ec6NV99KCWqmHAOFy8
6C0l7xsa80q6xTYhQUR/Wj3s0+z/IG/DE/mtFUsAMEII+lwIYCkeGdglXgemgpXe7yanvtLSY8C4
e2CpZL/OCMOCADjTFm5gfxXUs3cAa+0E87ScBBoyvvuSGwXz4zcmsfLkcB0LxV6T3g5BsoZmOTND
zqYY0vwjGpjsIy0iBknC6NTgZ59NpFDWUSmDLSg/uNgoRzetoD04PDVtxJudGs9BGaqPhwvJseP4
ErdeA6VenZR3vlavP+qLbcjKApDF07T3Jm8J78imn4CEsqs7y/CHtIibiVNTG4kXD2GrR1JWNl7E
N/AuTtA4kPHY0upCALP2m1y06wrW2tTPtSsHFQUkWBCVGfhqW9iWHfDfdIv9OKwvWhLEOsUmJ0sN
lV+6Plxm5vP5ZhlJxGnZVscYRPM5jkZwsO263hs+3HfDsfaMYKBI+ZxCP5erzKWE8wz60lCgKWTN
/9kum9FdPf6w8Jv1YZHNzmY4ZqGcSdMS+jNUP3EOo8oTsjWjzv8U52rqeV6udCsHvQbI58eS66oA
SuOz1zTTThxK0Wgz7xqHZjR210fVX4rI7NFWLkRURE7qQeHTk1X4cZXV3U6q+4VQ0Nxz+ZjnbT9G
uU9Hz0ZWg6pDA5rJeN2/q/7wofJIX1SDTrQcBjaG9L8mc5/1+ZbfJTKzaW76tOXYUcFHrxfnqcc8
HuD7UiY019mfcxMFUBgD4pHixmOEq9elNM8bXxaJfaW/XUbyUp7YCnBehumrep7vaAED3aA74Xwo
X1c9c5Ssld0+J+HpcrS/SHBL0cDolkgJwfUeZQtEqQe632GD0yI4asrruqvgBPZKi39SFk2enWN0
7dwCkRYVajSJHTaZEND8OTjnT7OJ3KzsbJSj6MIcQRuU9XnRKl+feXIvDjQwAzTFnkU0sldDU9sA
G57T5cJPNgPLSiumIJlMmPOlBbKbgQylbko+Yl6VJf0LMiQAfwO1HeL/82/GfR6R8a6TrCLZ5s1I
gweNqYQr7QUs2mTjYq7RkE5FRvDWDmGfzixP7wA6wFuJQpS1KxLb5RG2fbSv0nGjXj1kAT/z7sgV
c7GJLdbkqIQTAh8+C1/JVnIWylZWym6hxMtC+gPsJ73vvgxb7vwIAU78B54i57kyhlH5mYhDzg7K
Q3SzCXZIMt17lg6LfFhY2VlsGiDkvMYB7vJNftrZgCMHQh9upSbq3QmoYG0gK00ngWyOWM9AbfPj
OYCHb/ICLFzNJx5BmCW9rO/Zrlma01X46ANrlByiXFk/T93jY0equx9S/h7/tMQezbOn5epD+ki+
9pLnaIEcKF8h4Uv0xv7AFu7rp0qVFZjKSqqLgn48QR5OPmeIFeFxsWbyLt3Mh5KGFdsATJR/1YeE
sZwqHdV9TBNuuP31GYHrgUhU3YNpBrQ404mgiPGYnYoTEt0s+KyJFtlKN+7FxqEJmWMXy/+85gJu
TG7DHKUpRQb6Z2OAYxCB6Rs3YDZD4MC5VIsg0xlPCzaG8bPE5tRlzHSeiRg7Ug0tjtputnghCAXB
KecWOBCSeXHWNjQjyAXs29RGvEfZf3LI9DByGtjpsuVRkrJv00kYrQ1P7MICv0I6nDC3KJhjbnBb
VL3UEXG82zO6wHadIR9qNNmtxY60MCJlnJnRGCIePOwHqb/0AuxJQupjvLteLfeptCRWpiooNq3t
ik/AYXzWmH0be27PeGA1d5IOFn8c7vjeGUeHRqz+gKEFESh4zzrnb1H7PJkSHWUZiUwpnaBt3Qyp
xsmIRQ4o3BYEjccqN1dgQ04+KrIwQ54K4YxagEoSj4qjv1IeBh1ofdy/xwMqLgJFqP4OwgIAzPBT
6s/B+55CexU5e5pBPk2uDa16xifrppOZZoMPxHUjLpsLlXs+RGtbaU4S8FsdRjLHS/0UtxIPVOtp
WyGjNqVE9VJ5oyW0vFsU11de8G9qjFosSqzONCsGloasQYOM8ZLF+STaTIqLk2x0AmD00ZUMnc50
bK9WYVTsvVdjbADYDZJsI9vaYx9K0gDAiHIDlExCVOhpzB9z9DeiSTC3EOoVTCXFAoVVh+Rvk16T
RR0uCO6EoHdL/nV+DAsV3ONgNkFV2uomJzEaWOc5kM1EYEt7nT+QkYXImSkavmm4HhS7aPjjQ2aw
mgnURokLmx9IuDBQ++WMGq61vcQNNqXro6Npaf32/SFUO5S1GRkRr36xmhr/PU3WeRtXgbpiH3YI
Put0MeIXjY4Ku4o+5oXzA66Ana7xPEZcnKuUPf/8veMqHAXdgcVVxE0n/ZkzpypuV76TI6VQ/gsu
Pq53u+sjDBFJalZUGSrhre/j8/NZyJ5nx7fmkkpQK2LaoET1mBvTxHobalkIWiPS6+985HSdSwkh
rfJXqCAdfrBOv00JoxinbLVbEV8YHvcQ3F9meNODHUZOonFFM6pECmPb33xuW2qlfEB7z9/I6MZj
T5sKzcUjARCaO535jYV5iz7SN+UqCpKBNjVOy2om0Sw6zUuI3415ScIrsp624aK0qVJpbExv0DBG
fMVn2fvLvvt8Gb1GqhB7yEpEpNsQJvEwi2SeQ1Gy3HZf7J3OJt5Op7/mT40iOHMz8qwhv+oEqSrS
8Jd8K/Z+sgezEw7giwnooZyX8b+Ljlt4I7wMgmir+ovvB3J/Pu4FwQeEPI2CWuSr+EfQD3EzRBHx
e6+A5cCN3rhERMeyeltPU20ppM5ak20YT6XJPNHgHvKSFctMjp18dRJgP1qUumlGMgu3b8sZttfI
a8IdK9bItAD7Spp0fjV4ctUyH+GuL05tGmffOTjB4zTCjbEnJB+8PhapIer/a5xa5/Myllh/Io4J
MHGHB6bBAe8YI4mx0jAbNTF2ZzVnLaSykkyxCnvXfpFrn2ucB4P71B3Y1kWVn9vDKn3qkYFW8fw+
C6I0FnNOrMIy0o0+/pDZQzIVK3lyOo1L0Um+C6Ch/HaTTaOzsD/IAQ5ZVB81ELatvlNGQctpcWco
o2vBshOZhidMfZJDee9CLBcke03sBX5xczwdPkXUYAYyx9ett4e35iRmNpEDQhs8Oz1ObnWfhD39
u1l0SV9rJM8MHlMo6LL1fNPzafXFWXK5VzEdus4ejrLhMlDVYNUOOQ6S/EgCwBlm6qnI8d24OxC4
LiKUxsscybArx6U26b1r2jvtJNXgvHWpPPEXnAThh2BMiz2kn6UhzFIhEuF66xPLPpKllWplcZB4
kRhNJlw1SEOvOUpgKf2MbD5dPvD2uL4EDRa4T4iK3CB6SakO1jXnpg/QhFK3qkAgwXJvTZnVKpik
tBd1eYGuhRIGYMDxOgsmE762JabVesaJzxtKKgxIFbUFK2eDYOaF2b+KWgztNiNKk0ZTcb+0PxMX
slLnpqydMoT5VXbm18GDtkvSP51VO5SYaWuR922gG7f0Rr603mF2sGfo0q15+r3lF2LIenHBzBRj
frAV+qkiPs4ceBB4SJkzCwMGatd5kNI9Y3x812d9oCV0UX64EOgUt6k1gEMumKZuwxhCPFtHEOWk
1nEHKG1KXK7v9zWeCjkHxCMCQa87AW+W27DbAHxxxpkJiRMQoKCVy1Jpb4jtuP8Ox6+a7OcpHeIH
jLxjOgINXr710yloxpRLvRmCgLao1ByXah5lA4FfSATDa0vEIjVQiyq4x5m8aV8TCjEm5d5bGAxr
udPQUITUgyPphEp9iBXGN+xdO2cDxAF8UvI3FfO1jtICe07XQ1qn4JQGAbs3QCJUgtiUiyMmrBXc
KLXcykoGgYhhLYZUQbTQdyVRc0kGZtMlg+OyrGxoJ3zGPGLWEb8Djpdb4Pc08yr4OchnMIkEWG5R
FWBG+Thk++7X6fJKQZj1spFueIBm+1CaI3t3xC22xMB7eEWdtnCfPxEroukA0F7xbJNAQPEqYsgs
zanR0O75+j/yti6UZ53rkYOxHSik8wI1Cy5qFY1+g/w4qkbMs7in4/Daxx95hZLoEKuWPveKnN0R
nDgcQT4apOgcU9EJFCdMMmk1cOcQnHPTO940wuYWoINZnUmfRAOd9z2tcCTE0Jzv4CQAWnMLtB2I
Oj6vBbVBZQ+g2Q22tGNKdohTdKTGalxbFs7F5KTgmGproNavnSVk5rjM0XAsrG6Spn27Gz8LI+JK
VocyfDLZqVDCeAGCHdZEkbqtuWNdlpTVbnYKFHLyqbCkNcf1A0yB4OFwXYjeNerhMTwzWDvNRffD
w53Cy4ozUJNgNYsZ+lHFf2Ddb+7gNjU3VfBUzzWbV1RhfvZULoDwpyNDoOIsPfghcHCUV7zfpDyU
0ACiU/kkVnFziziuGuFdMUQrffDzWS8F1UmLDWNC5wikbTgp6J3qk+fYvh5ENHAvLItwGHt/SMrm
TiW1Xld3ljeHiGm7/2ap0abrxZQMcp/yZBCPKrvmZrlPuhxKEfM3mUpEhmUiQcSIRYEYZfW3Url1
Z9K1DhCTWB4I77FKUUg4Vq0vPBUpDhr5MI5NiwWHfT+n8GXr9zkq0VUToT1g99T52OTUARQ0B7XU
80gSNYSQpkJjf9BJnjGZA2D+egyi8rcOvD1NJE4TR5eYmM52q+4syBXswpJZRx8JXIh8TUx7qH3L
OdTKTxWLZKJ+nJGyyq5RWqvf6loJAdq/qfC1GufgNCey1OK4TS9rk4nZebfekc+sbx+FfUvWOlbs
opttmuPJQttqAdar3jpYwJaQsM1JYDmE95Rbqq6HoWPLqywTT6KnG02SZz7bgDcflo0dZhr9DbP6
Xs+QUgU4otMtgSqsT5jEeApZK1twLzbYuPjHjh4SUnNeE99tiUwiRk5KqWy/NUE1q2L1aVj0D7aS
B3KxxmoZXAR4RhnRnbHCe2cRwaIAvDkcqq8ptRdymZEqXpsQfhB4VqbylojIzPLyLjTGVvhamIu7
xgt/EhZeThMYeFDofgCHpyPADmBmaR9X1ArtQPbkcg5uYvpNLFAmMGvi4Rb4j/NMiDBo2b9rQ6HR
qSr5AWl/k7IcS0dbiqXjKgT87e9W/HydOIyBZ4pxNFRH8myJbqH9fFJHuaeCCxZEvBN9LEqSmRX1
/Y/80omTlgdGeNECJfaM2ij+RTTrcoIG6UDOnLGOnlnBbLraZ75KooqUZAQ2PMVDOXFzW4Zg3RJC
Wympzmdz4xjwsEjfK+Egz2VHyT3FueA1O+uE0WbpV1k0oYviJQx10aMRNExlUNkmH1Ks1SxAPYXj
mNorBmf0WmHEhEdCbRU6qUZdOvrmGwMJnJ41999FEsld80aRUGkZ0SITOcw1LYi8bliC0a+4mUmQ
tqpB7mSq4xGaOBF3IBzmcCgpv4DqoZvne3bBn+UI1EUOLz5ovlAiFrNNjDYVrhqGuYTmc0ev4QtI
s5/I3IQdUHdfQSMFVEG5NsXsNDZlT8rsQ/Xq5oKzmjIy87EXPcRQ6nTU9ZDAlpdrzs2/w0qmSEO0
cUVJduOcdsMofcMZ0LndNJ7LMNDzZuHivHphRqQEJE6LQkuf9xKbYnc+k0h99KXoRvTRrAZwrzo5
lEZj1xxN02zJ4QDPhGmoY4/ral1bobQs5Fi+toym9YeiiTtrEw43pq/cIcMYr2fiqDKQtgFpPUL6
h/NJlyQFtI1sPoKxHIErXLWvPDKMIGPVi3in1EsBaGkArmlm5FC10fTr57vQ0UaiMKyrWQ1FhigX
yklp7I4DuN6QrgQWiZrAIl2xRR7uSi2bCEL+tDHZDAtCwUcdji9WSTjs71WYPaiyEc0qs1toKcdW
gteeTlHM0WP21cyd/J2+TvxKg7US31lt7mnKmYBBasz8HtMJ3LUNkuzGH0kfiRlzfyo7tyOMFS26
IuqdU53Kdflptb6uGEUn7+XElnv3wLNa8Kv3e/rmZacdHOCpz9V5mlryX4pEZd2cQxsIbBRLWu08
2NYWSLeUv/1D9HyE+5jJEF8QDBjJ9ycHA3aXu6t4edx+TWZRtRBBOFCVFX52oTBYPmXL7+mNorfe
vk0sx12DRtHjrABJh360WeqfdlNFNpXxKJ/wPIQEoUW2QFmG82Rm+eGa7c1PQsFjevl7jvpCyg8C
ipt8YkxnsoEfDPt5UPnZhaB11HFgMxOichh/CLZ3N5GN2++0dh5s81MayJMizqy+EACSMgOWDE0l
DuFkwVw6sZQ610gKV0N1jFAJ7wVBMHxvB2mw2P2Cy64VPOorS2vvP5XtEtjLIfF8qLOm+YS3R0qo
fbLUIIVnurWYusHs2w0VNbtmBwLWjVKOjPhKcQ/1LbVzSFRoE52+DM42r+POQcXLzrPfYa+O1x6L
4Lek6ANjtvyaA2pJf9BlwFh1csze71KVKOwiJlSWzC3mBbl5SzSb/ZBQ2aTE8GsA/SQeQsCHciYL
PbGLRE5N77S2gC88275jjAcu47xMPcOkKIjghVE3tyiryY1zrl72+D7ucCvpQTDunfZ3oFi2VA2v
e7+QNz75nqhvEoveKW382g2oSyG5U71pCJETNuxA0oHUZtwC6KBRqZw9SJDi8iCZhMn50moAwDLE
Di+oi/DAoDY5047v1XWsMZc3649UfV42LWYX+6mNpHAQEYSo4SYm0i4/XkcSUZLMit9R0eygyH3/
j6ISViCRtcfb3nz+OZBddzUuD2gvHmJ0ZgDCo4bmcAAG7RMcnxh05sDmbuntNKGMNwGOOPzFP+J6
AvXx84rg6T6saqMJVqgMYAGF3ohvzPT8yO0MUksFGuH8qR6xeUIXQ4O3TVUagnNPG58mFnvl31jl
ndDIlwyKSc0WpHosQD9uZcr9li7VUb9hSVS7i05fvrd+wBZ3r+gJMAFA4g8ZC9Lon/ULNaoSrUE9
HikPUr3Eftkd+oMIMIkYU1NdB/ni/2tW0Vmva5gKw97ZWKkP804Zq2i2qTyVXTpbRJ2oI7k5B20H
G//ydNFV5KYyvcFg/yFM3dXmqFdlESh3j9e7g0npLjRBfzn85+EtP8eW1jZoxsqXksGfUkpYuiOr
dm0q2qXGM6ttoxPwytbDSEsa0l1uUuo+raFYt6lJ7ketNI36VAx0ecYBJKpOS5ekLBZsoQXE4TaG
1NRTWX/7zPkIKWpa34GVEIZKnUcBMuzT9a+APFPThBCCcHHDy1/0PSWljf1omhTrmpzwC+KmJmuo
v7/qNBje2ijrYhTX4UkVqupLE3uZO8IXiWUf9oBzYDeXQua9oXbjfP1LhCxLifcqtsPDFvKqniQS
SLtqarTpRD/2pCd09NoMCJbl5dMnNiNoW4zTbpPoDfHbuoV5H6NB5WWmJtnlGYnsHB5sFrPRcAXo
gDOsWco9O1Frg847apCHxCSmroF6fk9kvr+f7lKOSHP8OyT/uoXTr+2+2J4T96jiBqDNFbMEv2wS
Cs3xE2g69KCuNsrNuKPwSAveUsrftZwoVumPmP0tHY00eMw6lenZoMx4PpE2A5ckjuUev3Ga/96u
UI9cLZJO1kUvSuTgJa9SBrhZgv+yVgLftzvYLmg1OnA5259LsejkVit5gnNIBJLLex9lcUA7MOaN
aglfwvM0H5/l7QxsEY2UTNUtXc5X7vwHpkWHZb+zNncnm2vtXPRsmiCQS37AQTieb79L7fIkQn1R
5ztmWDzqnkHgnCy6JLUM1AKysl9wTSDLdXV5aybJo0m0CwdQNgcC4ZncN68+QKs/e5ojUfVALQPu
h4Jj4b1b4fbzUigvCuUWjsydNd2U1uIE/g/ck+RvZQ+m53sx2y0Pa1HZoidQtV8MK1R6akAKLmhR
srR1AuHTrIcSvxDQNgz2O8pSbuVxLUk8u2TJEBOnQ/R9E9a7enSv8m1OxIWQybsiSXqNstih3Awy
xpbdNqvN0UBH3clnRSodqPfIvDxik1wdwlLvzDWVWjFwpuK+9LnF/PEH5eXl08bAQCI/QSZceXui
hv3EkvCzGH9EPQp0rKG8aOGiWY2CZ3DTUuQz6lXUCKTu+W8uW9sJCXORcPjTdKhjmZFDw8rZzPJm
PGrPe4dQQUm0fz4tvQBtb4SVRiAljYXuAu64rGA/+HWENdgUqISJMsHGEmlGBG1XsFQDMBVBS9H6
GrOIBVSeLjYZqaiZ23XBSsNcTBbydAQfs58M85sVTyhrOVUMfATAmOIldAKQ6VZ/il890DVtedt5
0hnltpLE8W5PNPVe/LV1et3MgXF1/BxisGBM49bLg/MXa2b8cmiuhJmhSSeZbWCY4i1qQeZHH62m
AxZLT64sZEvrFAogMCvBaMKcdcIHWZNprfSPIN4Qo8pwhfkmx/oXEPj/MbmKHN87qv5Q7NevDcdk
SWvk9vq6lzsuHsfwjmPkn0pkH3IMemsJ+vVpombX+Z9X79xqQDnQD8+i/kX+PO+kCel5fnZdw7Cy
01aZTdd9PUgMUnPeImA3uHfeu3lbaDAfTp7fkxeR9HKpMAEEiUWIaSRVy4ahzqyC3xPTsTxoi7cn
B6VZmmAgMA2CEOz3ZLa6n2frQucUROTgixhPlNIpTDXyF0Z2GviDIxE4gnwKUYCHUXpHsDPr8CSa
EQaShbz7j7Ca5w8GnR6i560ElGMVyDnyWwxtRo3sUZcEvohbqnzZ6z+QpR7AQbZYfu4c+PskY3kW
HDd3OsxsDGo99bmFgIxvFF2jNndbnGwMMrxC4fCQdxNu9J17h6V6BBU4bmtDQhVL6ZnnFdOMAbJY
t6af9S3t1YNj5TuXOzz9CJv04u2ePKiBlhLR793Y8de6Savm8rxkRwxHdlt4WfgKm/R1IErI2zQy
LMziAF74zH0UuMJmZ0uQg4sh6osyY0hE9kg4XDdHd26xomVRDFz19OaJdkMgHWCnnJ9+R6DGRl2y
bm/70KkspMxen8MlqG1ly89FuELgkwtpe7BHVsPN8KpHS0UZ/aeW5MDu2yvanCv+UAo7V5pY0DPf
JUrn1zulUnLVEgqm7MlgP+Zy9mNRDR41JewsHBZc9bdbjjCg9lD39DIkK3L5Jsn+gNmfogtxuKk0
4yxVhS8HWu2TYtn5lTIWfrOqmJLetaYgoRC3usMmg3Z6FPZHZU7f3d3jYNGMZotE6DLv/B997+Pf
FRptzhFexHf8NLyhEdX9v8Xhr9X7/fuvZR/38RdPN5HtWe783NikcuUNgPa9X+HJcQ9v/WsLJqJ7
tumyMyPvaFxw8ksTeAYmMBUlJxrQ3uQSYhaLnlnkKtTUNa04SQ/+woHVG0lM0KmNAuAtkUXlSjCI
cQhA6gQsVoDa7p40L/sphhcu8IDk93bUHm8/rYs5wvyRK5SFsiNOpu7ybTFI3TG1AaQf8AIEV3wB
MAHBCuipLPsaynPYb4ROMTcUdIH7p5nw9kGLLgYgjXEZiM3w4UPIBYmg/qz9KSNvRRm5jauaAemr
kd4AiuD+Mb+a/Zk0GnkT+/Vmz+H1JZKKeeG5+0I9yiAeOWGeXC4EyOQauPkg1/ZVPn6YdEKYzt3l
kkUHfwFbgy3FDBKI3pb5nNaL6k/BeD2rhy8ZkQ5tHqHFf1SWJKAUONHtDWSU4EmlC9SEtaFv0BYN
JzLNAKkRHWgXXUG8jwZzNmm7Z+1GjOeszQ0XJBfCyy+Hu6Yny6iZ9trh4QrCsYnsbiAXdwJrOJXL
YvpbacBHA0t50CdhDORLn3fRz3H6/OvX/hiLWQu0EwFUvJjifj88+0QcxC+HpOuGUVeE4+e/lPZA
putkeP28zoBQ+JJkbvkAQjvGxr7yuYMAT7KgqkNcQbLb0crUwQwtyaOzOz2ftkycW01cxjsrh2pj
TwkGpnDINZqqgJuBaOUX4srftZsm/qRQPs64FErT70/0RYCNxAoEGQz/buS6e3KB539LGPpDZUi1
TqkvbrsOTvONsOW0eGZu6tSF4jC3xKqrXh5o/PoEuTvtxVC5lrig75dGE5kprGeLQQoPbFLSnH4y
AYelF6cWpWgyZK+1g1WXDTd1CKYjRO0iX7sg4VDMHzkY8kxadgNLb5o+VXjTP+hYCj4AAPgchHl7
A7KoXTEQQnH0iXmPdhCnZElTZBnbzSzeCLOz3TF/5jocTVmrHlKK6oUMi1EXN3Woj6KWRIep7bb7
HBJxGR1A34eqqX5WwwyDBV8jG4l1+WKRCakdViB4dkSYi5qkIoRiig0G6wgI4eHqYTzAsjIAFlyQ
P3RfNTslG1Dd/+Va+yfCadUZSLJFinLeiULku3OT0xw4awKgl41RLlcmIhm4lnyHz+FrBYMsSPhV
vJmNMk2srY9VPSEAKfid9OjAExJVarPbBfXieV813gxQX34lo9rWELjaRPvJ5o7sXZYuru3gIew2
RPhPYUQ/UCvqWxjAdxJhebqj2kX4Gjg4d844FnS6whC6I4jhw/dt512h6NSeAoRLPt4a9gsfTACy
zSJWv4uXobAvEMA8ONlWNL1C16LrXWMieTNJqIMSJL8R/ySIB0+lfnIWPw/pMU7osiX2EOlsGuzT
KmsJsvmx1F1c1067yF2SIWH/ccz5YaTCeIbh3VV1VP3ZNbonb1xnGpZYVkOpLChwF+gAuQo+X8KS
c1FuSMcwP88x4e8hMSHkc5Zg6U0L9WnfW+YYH65/zXdz9awjNW/htwhxAdEHcew9ClsgaSfyi555
UKgeS7unFR+m7K1YbhHwabLWkQvk5E+rLleocoxni6rxNIUipBUxg3UIzNLaqnzjR4ARLMwnUHfV
cPgS4U/E8JOE9mA2fk/Ko7X5v7h+qutJka9Ng59aV969kMngNZUoO0SGrD4hPIb2TyKpBlPYFEb9
8jBjYnjfIPjXq/e4azA+jpcole9WpK44aPkHmAQnjL1f4tfm8IrpiLzXKebR0G3wD3ig4r6WPYvu
ZG37VG3TlfCjYgCzhA0vxYe+08oiQPccDGLpeEinB082DDR71amMTJI7D12hy2DmjhS6F5aY52aA
R5i6oR19mZZovKneIEj43bDZAnPsQjkG93XaTMJCK9Wm2Q+FSEadOtcc01oyjYeArdSZDPQDPiwU
UYSXiUJEvujTo9/YcebkRqt7s0+IDU0ysqwJsdGcIpjEn+AuzeGf52ZNZh/uy9mrDXO57dDRwqw+
5zC46u+/gGqj5AofMxW9HKyfwy1ac7iv2ufOab/XUKr10yT6Bs12r//bzh7Aw4BLyOli3LLGR7YN
8cIRU6YemexNH25SVdL2p09xHXoPAN7NaEHg/CtqD+kf+mH4wEKWBXZT/J8tq/sWvWq1p8WKmeWd
l7y7E5DI8DwwWFE6UPnu0O7+w4M2J1chvVrAi72Saan/M2AzUJdveZS6+dzE4AkblNHZUUx7cJx4
9JokM/mA1/R/Y03RbTW/8msYNfy+q/j1ySRxxxdyKucgzTitLHFri1Y79W/SSHKIH8ycf+pt1W6U
6VQ+BXIbVVHvV7TPV5ktuAX+pgpgVS4IXgQVIJz1/nLL0Nxz64hnzTyzJemJ/0RGIMyg3yFuzMjr
QZTAatpJfubaSLrmjEht3wUMQg4j3fDVcyA2kpwrN6bwanEo/2l1SZrLNRFeBEQJR9e6xgvkYpsX
5lSQ4fMoM9sJHGq5mhmvTdlUAGPUPdn+szgkwRo8DvhDlgyWnBIrB3/uCRYnHX0jQGeYCweiCFrP
9dsO6CYuZZTudJqxgut8A+7LvJz37okH+oAW7ajV3h0RG6YJF9LncGEpH+9kz21cUFScrGKqgA78
KtGVF3SLDSWcLuF78MaUusQjhKH4CY6RWTnNVY4FK/NXYQYT4tJxLJdlgKzkne0+pLiR1aJ8ZPH+
Uc7H1+JyF/3EQoF/L8Z/l45ZN2GezPqek6/ZZtw20JApUGaQF/I8TV9R/3nTf3kPSnl5IiTOvygp
XqmXpMQeuvwEsZqFiSztxn1wsSC5ncW99V/20B/2e/d9w1K1dC4872rSsnQCZ+44ZjWzBxjTu7we
uATly9vKEcOutYf4C4ZvlB59drFAEwstB9C0PjnhVsLArnKJtkBRME8OYGAMjFxv7tsK9tT760Rj
nXzlNQS6SuepeknoaFFttZlzokAQoowlKG8k36PUx12K68rjzRK+0MZTezt9Sha8JTzpIKKiVWZq
QjxAx6UFxPqs6SHz5laz5iuiM/XlRJgyxYkGkfjQLxreEBqYJL0ssvc+S/O89k7NDJ936RAPHT7c
GT2dCfyuJxSL7YJ0vozrtE1aj4wZbQg2mKzJbUzBD6PGsIZCS6nAPMf7D2Gj3S1VMRyIYvrK3ki/
vCuUwtFbYIYB+v74o+uVya2LCsGXfWuNXeof9TgpHUaynDUE+YS/Oy87eNueEpeUj4ezzJx5EGXY
43a5PSWEuc5xSIp9kB5JvfYhVuokq67sHC9KzO9P0vKulFeyk9K1Az532AimIvoUPfQxi+P1sujC
CRf2+zzuSH4Ocjrl+pisNPfcBeiGB0nxdmaXhH0HZUVyJBqJ44q7ZsRiN+6bin7Tvvz48WYpgSMD
Y5ew6fGfcMd6roU0FhUaVcdqKOVu1kvUsUWXInslPd9N4WoPhsTJSSjDlraftjJNHUlnlvcISf/c
Q8888IaFx+OSl8gGRpD9oaRyEfo1UU0/jEOiriZsHdOBNgQew0cwjyAJVcpxXLBCMpyjYx2AwdWd
ETds1vkd3tcWmg3Qoy0S3nw6iPMPIUxGNkDpFFtBP+GwuZuLORZ7DoxvrsqvuAu+marMuempA3xH
V0BSjwY/vJX6xfQ8rPaFA3deHwGIOKaKxwlO7LhOTO9U3zHf5d9llSTLJqUo4jUhWOaX4AEfM1U3
zuL3fLx8VgHW806Xlhr+mLKYS/4RYRvfyRIN8FLOnYxrKm0x5NnskIhHL59mty3EwO4BB42US2oL
bZ7UncOcG1Pni+hTWBnqnd96JUkRaBmto/g8eYiVilpcQvK14fbI/8nbf1KO95bTB+FaNPCs6rcW
LVzbwvGIU7AYSvOqfAaJj5WsX7bX17VxzNdpEjm0+caJl7AS3TQ/9b6XDAXSTn/cG1AEN9Lh7QjV
x+t6cieIqwJR429W5kwm+c/bVcAYWhftzu/rkedjbJuo8rkWUu8lbKNhdpFweDN4iTpk7FHbwRwx
fofE/kBf5CzepjOYNCDGNGuTGyKROR5ZzAgsD0O7sZGzLxTy2+BfHKnbjI7Rmxvz7TpuXF/k5h4r
vx+1wfLtj5OV4UpzxHY+ODPNXOW++FN2gAJVvbaenipIi6Aw/RnN+ODm1U4TqdqruG+4SnZ0PMBB
/dFkNLtKJqMWw9DMuzbrh8rdOq2B7gFh7xC7TmrIhHCyDckakhenjuX2T3StW+DYY4F7q42MHlMR
k9w8+Pt9o3hXnu7zhiPGrUahslI53ROiJs9+zGJqd2Cc1yNtB0LQ9HGSC1PVo82RnBxE4t2X5wYw
Ka+aAS6Odtt0L3PYXVOZJgUSZIML+wFVtZqzFLpX62Ejz/+Ft2T/mfeOHZW/IZJCdm0jjLnGZoKg
EFBf8qChKp5AmWw472WvYjDuTuNq9psFR1dtK4XJmatwxyPsDF8dCIZIey6QLLfZgCorbBYEOkd2
BUZSX6e6KU+HmFPofqBm4g/NCkbL73E3ZNYwbzKEaXqwJQeH7wiGQ4jLymMOy/+3InQxoZkhQz8P
o/LP+vQ3pmN+gG2JqkXWOzZnS7s22isftXCyyHt4KIKnsI1hy1MoXGjAuL8zNynXqiodp+EUs8c/
NQco7wkivgEgSs+8LD0Oxko7IKjuLrfF3ZL5CCPrZTlvdw5dDQmP4wKuq8BJbxf8LgtgBsi1j8nO
qVkPmCr4hFAT/EptFQ3Qm6VdbQe/8dyjDW+bQJR5+NgUS/GPZoJD5LJ3aYBJd1ScYRhLQwHnAEGI
G5jk4SAPj74SN/Q+5fJlvYNJeuMl5hup3GAfYs6wdlp1JBoPHAHHhVOfQTPq9Sh/E825ByahMtwX
lh1M6TsxRpWzmukg5OLgaBTi1IyM/iOf4nb5N/rdi8VLlQDY2yO58KIyo23jsAOLT0U699ck2Q+W
b1C/QgbeK/mpwoi2VF4PE2gy36N868W4jET+XXF93mn4HizC7CmEbcRacoH5cvPgdZjXyhGZSQv0
0gdnNAs2exazAG2PRKIOzAdrVuCpdVgXbGRFmbWjBWZzPME9idy7o/H883Vjd8qpBm1Mg34JRwgZ
eUy+O1jWO/59EkpzSjLBdofNYP2lguKKr8REFTJB+uzhXkuW1WSqQNUI3SM66AzO4gPI+sZiKIHH
7xJp37WA8ksNB7ofL0Nl1cjj8uBTmwdcMi/jwLbsWAipmMxswSQ1EpF1CJNWqk95C0/S0DKSKeS9
AajuC6AzooUY10O/kRJw1TnF6qcFR/ZvFORBWc8m0/cSqcDg99j9leA9LX+lac/LaagmQ54AIJw7
qd17Er6fW53ucwkva3RPHyRWDCSD5JqiIfDbCVovC+4EqnZVaLv5pkVSH4Icq4dZZpc8DUymXl8o
92aqnxGGzrl6dmT3DhqeYKOCkFzuMAJLBXeNQL3zl/uO8E6+LJ9x90S68kKTC8DeCBekf3ajhs4x
gADWY02hTSzq9MUbm9D16HUw1B+rH3ybnDik4UmyD6+lsS6j5EUeCQYPY6udOmPmJFkTRdeWS46v
ET4yi8as2O8E4A+1peu3qEb9Jg2kMznh5VubIeNVsMArY3pogMhdU8A93bC4NuYE5i5NL/ztL5UY
Za7FT42VYvrQTpLaMVGy/LLx0ZePCbv6nSDtgk5VBnMk31+hRL9ALDjMDaVvZWwEl+QoL28977d2
kTuL9dvTnbsvPE39SHlNAIdzkxCSex5kiT8rZ7urAM7RYA6W9TqcYsYVMbTI9ewCp5QBTCqUQS0a
9/I5YPJ89vtlj1Otm78MrTz7Us3ap9QMg75slZjaC/HXr5ajPj49X+ZX+7bN+aKDOhzTm2OjxZ/M
bqv4jwwuv0qKqcyKeaiqLwQh6zSk2UXl8rT/azoVY6RKNNn2IYxV03mCMVIjn4Z6mlryUV3rpka6
O6eVHUMBJu13uDokPeyhyzc6Rzrnz5Q632Rb8C8JXkK73ju/rlD/+0jx9uRj2JDxemdOZOyTievE
DJMph6xygs4ZQDiDI7zRczsZE0YgWWiK02YseqkGLKZjF/qgXKyctEW4ydnc3wuHBMTyZ8muv27d
HX/nZMjTGuJlLrt+Nij8FdHBkdDQHFYeDUyPZlYILcd5lLSII8hGK9VuhsO8o3zHTnpVPQNqp0TE
ZPVxZnsa1uAWfKs8iHccblPDbSKcmkYo5ligPRhFLDt3KWILrBIZrJA72Gn55GAwPly0ryJs3mni
UwDHKs8b1WfoZXRzlAcBA25BOC1JcOSIv7lOsfCQI6cCmAZl7KkE3xCcbnU/rplzFeRo40yMhZyF
Z3rBRwNeJLVDx0AL7VvodswUOJEZWCfc7B7sXFwXV8EwaTGGcd14nUV+K7mT/LtIllY+F0MjZnSR
maIZLvHG3QD+IH6u3Oal5A722MpMZSqQc+bPecuoWrHP3p/tu1yKn1A4nQzTAivxrbarKWr0aZuo
XNxSa3NU4XVMb37NCy/GhkB/EsRf8Ljh8xd9gPlRaJ5451pBB7RKZb4PqDF9cc6IU5YDDJUg+TTW
+TzJm+Dr01DCpQA5+Ar6KMmFbvaDOHvGHQ/v1frI9rN300dn5I9ZrcwdCJUVGNz+Bfunq6DlqKAL
RJBjlarYEPSWFB257d8agMm9ns6sIJjOVAFNwPZVI3VdkBpFktbJQnvsv67m9j5AMO8xCwrBmBG+
mpx22SJ/PVzYKCYZkPwQweYC/tSQzTtVZiPlABPJms0lbW2aqzI9fzPZutu4+bgUS8s2mnai5ueP
+cJuv0Dbl+UpWetfdXMZT2mddO7SYAJxlJd+EO85o9p6pjclYnbbwEyi73e3nONBJqL7hyNd66IX
4ImGYR992GLrG20DJ8ojByVTWGYQLr6gin3mI4fHeJCTxxbmbrDVQaa7m8h2gWbR6qUj25is48Dk
kGisaIeFifkyRypKFiIoWjDtQFS3EwB9ipYFO9PXcc20g3oiVPpfgLFAazgT8vC70EBZtJbiBzKA
KzpMdAoU6WqGa1/b2iHCh2l2PoOFsaocj2Mkla+fqVjeqyH+6IJvpEfPUItJcxM23a9n7r6vXD3C
Il2TbpEDlYHHxri+JR+7lbjM20njkquVUT01F+sQpTYOcsAQctzN8TcSnGU9UQQfvXznfDNb2kJd
4AUttvYpE4ABj2U86YPBP1gog5n81vzqPrt0nRt9pKV1oS2MY5fadUSlCdhzdkjfs38WI0ROH5aX
VZBgdRqnpCnPgomWsD7jIIscHv7PkH1ECEsuuDIpz5KEPToGPTUxyB6k0na4lZhpruQKOPiMCi2i
fWGY7mHFPrnAvSvfa8uc7dLedVWaDjUrE1K9LA/u5B07Il78qzUIqeW5kQLMf9uJSF2aqeyE4fof
Hgc1T2RYbtzPh8uPq26v7WLlITlOzhurmewE1tsRs4NtGTdsbwnGCHQvQ2wvfLNmSA8I0qEGS49q
cdeuNM4om4kNjbA4yzZASvJWzQkI+uofYnEyat+VhEYTYLb9FsqEGRai5HTrLDC2k/v7SJFc/DW0
jbC5loz+1bmyfwJC1k6ig4HEyvtaQZbDR+4utEi22Cp2yMvvkJXhgNig3fUbTYn/6tTjGZlQLaCa
We4479X5UHtmELtRCJOcFIKCOOy8u3skUYjdUpajJnWWPwh1hMvhsS+gs9US2dkwqNhAJhWrgGTW
O+T25dVGOOKFetom6R4mux0cHwCyyaOsLrEGX9XVlqBE6xJB94MjL4w6jdiD2XPX84op4/Go74tA
XssmN3cpN4nIpHQXsQtfxoHOz8eNZpMgWCbfj11/RkbxcwqQ4kuvRo5gv9CgE8dhlXuVymSZyf87
e7tizxo23MNPKTLf5vsh2HuyI1SQ1cYvGr02pQx6RFR8UDLB4BJDAfPdqlN81GjzcaUgTfb4LH/g
03O7OvNAS0OkJAlqlDAwjfrbJ6WNH9JRWJ70qtgCv1h8EPB8qfqLKyEyf+vSW/kfHHm9UE9btXed
IG4G3MypQGHylUiXjS2MtIjA6zMnL5mUEx9B5pGdjpMBYbBvOVKSLJge8hZFfO+Lhx2RYdTKZZje
sYAOiFOGq7Rs2v7/Wqp/lzG3xXYhe2HQO7ILUg1lrXkDSuv4rkU6BK5cfrs0SURfaAMqXIfBFNi3
NBl99DWZoYo1t0Fpm/0DVpZCaWLBRoEK6jpEbqg0M+p45dk89QBoxaCRJ9LzNVvk4oyegYYU/8Bf
7tFXaG01eBlq838+2vW3xLsr6ZW71p5v8pMVW7NzVsGBTtRINfF7yyoGcp4MjJktQExQrgIaZfwC
8xVrBNvMVOl2u1u+e8L3A2so5KVReqIi9RWZdKvYJUw8gy3fTpksgkD9m7WbWe7L/I9aTmygsIC/
4ZXCQ+LjPFENSw1tZXLZINNNicPC6paIZxpFPGg6de9uxXNGE4KFXbZWv/PuJD6UCZngwpXiDFnD
cRuhGZRuGAaBUn0Q83jsW1I2ZGLNnStgKgxIFt173TTLFjOQD1rZSe/xUs/Sd3k+cHn8Ah3xWkvq
QNlT7sD5Hi4+WKSJRAwXrsOjRjNKkJMdRcX+W5268r0YM4MfO+4IM7GG1hVgqVPS+JF9yjBY0guJ
Wce+vKiROYocwR9pdrdU8MlPbcgscM3bdUy4A/qjuyF8R96Glfp4ZSuGhbXRqzTKqutl0egIMOXW
zh3YCqnCxVcUEwJ7Q70dwLWGQTAweXg2mOti5rePS9RzLb9t/5z+1EWvwssX6ctCtWhB1npclMTy
DBhw43sdBpNUh0/75g2wUEpBjoS2q7vdfqzoWaK2VzGNVX5nPuppBVYjirLBQkVcJiiTywqLbe54
r2uvI2BLrYQCok8jB4XgqSxE+1POa4FU0i3kx5Q+AQGdkwP5Eu+I/p4A5VecmHM0s0QVhks5GXUo
sMeRabNxSNKvLoCuKt6g36FUguxkPDwnmwQvu697nz31dvxftPNWodi8Ec4ZCm6ykPzqt2Kt+5Bz
l/5KatMvmBEbWX9ksBl+309CBK5CZFNGU0kAHZHCclv1Yha7gHtUQF7qwKmBgA4su4zB0sYRoTps
wgnP/jhEUOBGbdkqo3kspRBkPqy0v8tCClsjnHmrs6KW/w9AWg91og32Syl1pJfcuE0mNPNlwUEV
6gj5uxGLzyS4sD3TOp3VimU17jsCQplKa3j0ODtIBJP62chArwLQH8kZNCP8mMcVXlHPpwYc6fRk
3/dt2nTVkDEBMOfqK55VFva70bnTiUcQWPZEzYugQksPC1MbkQrZ9r1+73fSBfKNcZof4KgbNhwQ
u0yJ6WzuPx9UyaOZdxfeaHFVp26WAh5hcFRwz8g1W2gTEsHT/8+cQoKTaSMJBgwSlYdPgVu2h+Rc
BdsZH0FGCgnlQlYySD68IfgMOozDFQ0c/6LmS20Pg97ZwcNVvOL+pC5B0EF/XIOJXfAbPqRxvrce
hCRAmHYyXiTGZRMEdmwHPkP/JH58VKwaEoaYYVme+aeI1jutvlF2NR+WwsLd5q/SnyGtfr1qIbEW
ZzYw6D2MDQSEXhDLBZ0bOO5jejqjCZX9TLoY4Qxn5T5FYun81VGDyLFaCl3oH03M1/CMYbqGyhgx
W38qQJgPY0d+CDC3qS6g3QzukaTOvKBSSKhZW4rhY6aX5KonzS3WArURKmn2WMq46aVlA/B99bf5
aSN1qrzZkfom18wuD4XRI21Ne4XBM1Ya0Kci2l1eFEhdowckbA+sxzjzvlL8BAraimb+7O2JmuvM
2SxTi2k8ek/0bvGjgwN9D9b6/fwVJlNyt/gGeeSiR8iKHdYpe+WQJqZDYzZjGBGthcid2ZLr+CdX
6sxb3vmPiZwUMtAcpVFbCbjEVFnzyrJJdKNWM7MHlGDf9lZKcK8YGbMwQYjiI/aAk2IEk1KribOK
GEM/Db2PXArilcJlFFp2zOGe6/rmWqN8GHmycoiJWN8F8oel7xRqEDd4Lp/AmbRzfIqpkFKYCijz
LfHammEmSFUCi8ivblKUvtt8Y6gNXuveO6AMbaiS+KDkxamf17IGVwRXF2X9Z7O+8NIIxlAYsIqC
1daCpygvz0BfuBvqt8nG/H9mvS9kBWtkjhhowepYuZpnUU79mLsUwZaRRaBBBNuZVKVYIuf80/Of
g07MlL/Btd5rIWvWcXwv2qZt9bBbBkNATdQPQ2ni9ZKV3+nbcWN8xM3kCIUGtGZmki/6bW3IVbx5
aAB/60CwnmEIIGFsvlPcyfjjqQRQokcq2QcWGhPV2lJ/hqBetM0JOaaL9YpvMSt8YnaArro97FId
IxcTNsXqFj4ClYwt0QusyxPBnJlKqhNicK6shnEHTMKf7lQHT50HEDbDw9zRXWTRhJZg4M+dug9i
+F7g9j5SY0jDyHJgu94MFo5LjLeKVShxuPtRpWVpqfsBEGuOQl6eZDiaUzgV68I0G0NWlit+pZRJ
ilrkahulsZcjHOUOa/ZYC8Ya6X9PLBlEzFyX5XDYh/+MAxGND4o5+pFyndpSsv0T0HP/PXzCUv2B
gS/q0r2KtYyKuV7DTZavrI8E6+8DCgZt5WUlsCW5dnD/n05wD6oyU7UwNXNOwHGMfJwH6NSiSHLR
JKsa47+xPmjoovEtjxHt9fjV98T1ZSWlMgObuPT5AszDagh5JgF6gDAH3zyJz3KfKdTHQNWKSPy0
OC9PU4/w1jMC+L6zY/zDy5aqSOG0BQgNPN5WIglIEPSeCTW+FaorC/qykecE72RlfTnSa6t8HU7Q
OuWJd48cSCCzSXAst/NRa0+tCzfAZIwT4pd4duWsrmtcUhy2h1msuwIhpcu1g/l98zYSxSvG8ya9
GntDl12JOxH5u4n4GbgvjrvfxZVpGBLZ6uP3FFvTA9jVA7sRNoxXmDA+BdVCvNgfxLXxGmfete3T
nhHg9yGZD84/QbaAdQQAKA7o1eQ9/lany19ggov2YzRBcMFO6SceL4MdJq79hQifR9pu3ey+uiZz
HjOvMrYri+oLXLKR4xPA7qu/C2k0ZjlgDuuGbFs0h6RbLLw0tmC6N22GAB1kBRJbI4GbWXj5cdqO
AdvqANqIlYFwNsBivCrcRjkYWUxOZbx1yeA9KHs9DG3zItlwCLD77oAhKU07zV2x+vPw7utch2ai
CFSo3qtQ+iGwLizO9ZsenOr5ryv4thqmOQh2OW85jnXw1kJoD/JD6ivu9HFX0/riIXXK1RLmWej1
9U0Fm+StztekWcGuBwpooVvzEqabGdAkfyUZ0uOMW7UwIPhtZUSf7XPGzt0YkgZ1lRabdRHOKHv3
NcrLGDZS1kLAN7jEgR5fznR3s0sI5/4DrhQGBMi1puX42o5+4gxJ7l7twp34sLcXwqHZ1SBwLdpH
HnanHCPsAvDilOuQgcTAFKczsmjeET4pBurEVHkcu2DW8IHVJD1Vnhue2E7jbKXjHYHboUwimPFU
OP97fGmqP5Uynv7iP8O66bQUVK8WFswzSSZTuFoIpmTxgynEYInuROiutAIY+AH9MaBXqmLZ7iHy
evGjgfFzr0Hj9gU/E7DYdtZ6dtK4Cuq68cLKjxhrLS1Zn9JmRvaEiusnopO/pS1AqVFtlpLbRw81
Jz4S/n2jMWPWtG7I7rHQSsPOZKWk7pSZcVOxMVguIMieSA24op4Bycq/EEAABIyumDsrtkYRzvsm
Be58/DUmuUQqF542dzLmkiES8IRqj3/D2euKAx56bAL+/wez/+7FCLsMbwoGEG4OAzmOCccZAPkr
uD7f2zrVwsacdWmBPoRGcFnDxTq/gTruthBLiOUA2ictLGrRMw+T2LQxIIddQugFW5y8GX3T8fwA
KMbBLJXXreKTEEHYjf/PZz4WRaIXvnev18q+faKg3E44aYY6F8B9LWbjcaq7kwk+RQhHkV/5842M
MW3sUzPWe0DPQSoXPfZ+vP/5HbTWCDDQ+wtDZPOBgoMznkNvdP3cyfKWRGFc7aPdqCKF1NvgN862
vLM/+ILPE6vP8XZTEA+Y7KIgpMN0bfgei6VeByC0b5WSEzDPsCyKXhq5pitIAu2BiAENQMbrKWXR
NSKQ9dVWpMkKDB7Ek317gch2VS3eG2Qv8ffZcB2XaIqlrmbcz+ChNCTvgx8kecB5FbzE38HChWiz
oVNA7jht0VSZ/c3YiInN3gA1ld0o09dsHE2/DHyB7UQnxi4A2ki2l/lKBKjcguNCzILFaJqk3o/m
EMV1A9AR18KmObh4oW11BOktGO+0BCqD5IsWvUHT9Kn9lN00HKS+efjPgJwu5x53xuDfmaqS0rkd
gsfGlfwpHBloB+8fD4mS/6WzljcyP+d0RfPy7SzCHiwwlveRn/OzdOVAgKZnJww2yuKzMJb6b59E
2DTHx0k9gLePbXVQ6xeEdFCzJfzekvB5T8mmHWuMWLEcOkg5NiWLuxil1aOy32WaThubsPjUWgXO
mIkMbvQDV+TCjW0e2rV8+E1q85xjZAZ8/EQj8rV2746oDtn4D2QjkvfqxCA7hri8fbi0MIEGzvPQ
bOl/CfvMpuuCmunmgnaqv+BztRbpqw+Wa1q6VNsnpJCl4c0Au6poAZNR23KfsSqq1uN/d6eVp+k+
gf6vF0du3Rc1LLF1qYIfEIOjuqT0WKzeDrnMyCy/4LwVn/NH9uuaZylWNd6AUZjezBfiX0TOOiF/
vZcYRWFLwkV7zXSl+fJWyA5U2eH/BFLT199A/KD9jLOD8iXu6kPOxfStdFu6iF3iG0DWumRgZXI/
YjA+eH0iZoZ8NpNiU0/cFPUHWCcM2AjQsdIfgNxJuH+fEuu4ClOO9YU/cIjDQ9L176vLFtTQR2W+
QMhWmVumNIrdu+k7wGGGw++4VWtnrR8l5eoHldOC02Wq6fFwsXA/darzbalkOlFBbtwxXIBnwT1o
RTrdn5n+TcPXNhlIdCzvuPP01+AzFxz/8eRbgIp0dADzP0FD+E0ixfhtN1EbzQkl/7JQybFrblj4
aCAj5fMNp1rc7yA9+53QOY5js4teJxo2oSrjGC+QnXfjU1aIb70irtB5Y9JljKxiXLRaSaY000DB
xbcYgJ3RpA3la/Bw0XPL1o71Bo0fr8nqkaENaIG9Pl/YKb9DDZStdjEYuhMx97usjglekP9jCsYI
4NnKZXHSXrnOPFdvfQl1IJ4VEIY/VtI5ZmiA+A21SK7sZzkHY43GUUSlPAHm7KZFjKNsF6q4YOJQ
dgGVn8Rk/Jq43mD7IFNGjntRUXgdRyLl87SZ3i5vLWNwayUmQkD8K/FFoPPh8PJkrs+Yu1u8OiDx
QjDq+o9AV2HZCfFW2CW7iYWxMduR4vzu5A4p8wQXrIQQyd3jGo8hvGZKxsJudr8KXci/sExc2bIa
L7sil+poHt3Fgf/R0LFzbhxykxEJp5rvS87RHTeufRsSIJmScr76V9FV6/YrU4uDh6+aX2nVjkMU
DpVk1p9P/UusgWeq4twaIJ0yz0q0Wktz2acPWxV/uUIdxNciEBYoMQOZzML6azhJWTy95rKSimAE
2S4LgX82dy4TFCcsa7sh78Jug45324RIO5q3OTmJC0hJH1OKd/yea8NupdIo4+pcmv7RaPBgIe+d
cMeATf/Yljjr5Y86pJv5JgX65hECy0FUQgE0F8sKuyzlPB8+eCQRCFdpXByOVjD0q40BYTs28Wn5
ubT6trcTW41xO2Zq5k44EsvGbIFLpAH0gEi+jJxTxw4oMXI/W/wpvTn5f1IS4Ptg5+KeWRWz2Uog
JTGCLPZwoE9LA1Dk8p1he8Lx25ChyMsan6LOUf052JQpeoeD/FQt10eYIVxC6dQSg2bhPDTfofqB
GYppaiokl/U0WxMSSzlt/j9bwgJr/KsikDRJgtHc0PCeqhqy7k9pWhzgT0Kv+J7wPgw6z+gFkGoM
b3Aq5kTXysxLU17c2XvnfYh+20NMPEyuISfL0MXVgdJdStaGYBaCgnoPO5gxEKaReNMiStOWXuUB
pgu48jvTIpYG/wI4tm7/AY7WbIvZ+IyDMKnMFWXGyK0qEyMALpIYBZs653/RX5FldGDsLbS/FVS9
KNoZVzACnr4KuPisTmXkGHZQorz8yVV/C1OShy66cz/LRtoYA1ZIeO7x1dvlPqJFxJYf37SukjVM
KyKkcLi3r2eYmf/dEzG4T1HFIoarw9QTG9U1/1bIstKGPN0lkuecqmz/cXODVd0ZPhKh1NjRmaWw
mWElOKLkXqmtvpPvRt7K1U6hgYwolcLfGCLQlwVxeZjFokUJlUR5N485Flx3F44Dfg+MQR/TD8vX
GXtpfxVYMaS3dSzCJsf1/G3I1pmWH3oDPWX02j2TCX77BWLH1Up3pvq7t35SeKi5FIR38pXLiYYJ
b5e1otemu5nRyeomfl8R782SSSjfVr4V+0QXtuhg42P0mLKhj2EU5nZs5GXBc5r6BTY8wJeStQ9Y
Dnik1dEcMvtijdTCVZFCmC9rQ+63rf/pNekG73zjMk9GxqJvOAqFVIa8I4SxNtnY0obAS/4RoWmv
IxunJfp5QvquVZ6VuuCx4eshuyPKStc7tk8oPao5CDvM7AOG+KwXywLDl9daoRutw4vHVvjTckDj
3XY1zO44wkRtuKy0PgGf9AbPgFyMVRoNEabfzBa354uvRPu2JNWXT7XFW8TsRKDPYPj8EsHp5jPX
arNhGMnwBs7k9jcmZx9lBWTxyDkWdZZtkIlp6/aRH1dxAd5W+zVFzpBIA5F57tOicAmOM2sGGak+
a2bHLCQl805CWRWs3hRmRjIcEKOK6Xb2KmWn7EEc/AE5v9u2AMJEYdwYMFobJCllTOFIy6TCzP2A
mwONZs2k9K3CG4Neqwbid3aVqkkJUpkkChzNrFqHMCSwPnccc2aDc7BW2wHWnnQAnD4wR3E3gd+B
IzyTRUVJky0+J7GP5wMU8Oc8p8s8/8PpnllvGZknmXeiJ0pyimhTPZ+ACJvkBMqAFvJJ+fQXZj2n
gPEARBlLBHQc/vIN+oEzg6oOU6j8MO3mMVFaLn3OcnQHt+GwwM2CmiHitMJvmjFftkNKh9qRLQU5
qLCDG2tmU+5lxqvJd05f7PtNfNfIy7A/D9qL8cg0UTquQ4LNNLHp4wzNRGOkfnKr0WzPQplficMs
T2pVJch4sN/ZJ/yLz9UqJdgxYoGYBdi5ABwSg5mV4+SQ5Ow7xbfgDPAbqDUdovB8RcIrI9IUdkai
HYAcVrZFO1rOjfP/LnLmpLdo1VcFv28edoG//YxM66rdT4omjZ0JyorJHWDBF4QIBMfEEqDVJaam
mbbU1N/3Sy9crGrV6M6aomaTfHkZxIp5FLWsMS8rbKiGLCNGvDOVndYLtdF9qlPY5cBdn9f4Q0iB
Q6e3Hhh9cIuc58r+AevmSQGHwyPItADLzabO6TrSw59T9gWsjtWRls7sz05/EsGiZTxpD9/Em+pw
mefJhdU8uSimn70emGEUcy8fg1nrqC7XVviFhzLh6Q2zpqKHt1PItSORiz2WdX8YJ+11rY+xcnNr
ZlwMMvMEtClQ5evT+HFSj4qA/M6/u83MMnasnHqHlRkoFTY9K/mm9UV95EqLG0jb7SYLE4H94piz
C/150RUU3Sk7+P1868Hu89qZoDv9xzxaN0m2THEb7lXwkMlrWn5kArqq1s/yevTrFWPZsmE70TXd
xlT0I3Br1GQwecOnuc9pqoBezXS0mT2UUUDbXZdII8gh6BY4cLXxJI62Km7qRRL+CIC+WNHz8cPB
x6u3s1MFTXsboQNzF+1g4DZfnY01u1BWt9I1x9OU8j4tsFbsjQLowkjw6NIMOyDK+VowyaQVMqFn
O/dy3eQ3vHfoQz7aLeiz0qCQsfrEBhu1P+DuMSqRXp0BSJ2N2BX7qRxbOnGYNbDhInOnFmBOw+wQ
T4w0Z4ptwnakQBDpFDMUHXgPPsnd18lUeFjGYsmmCzNogL4pn3O36aOqlEOk5vXTo56YUlGmSZb7
yzSuvprYB8stZqtRsBMtt4+6+lGAfSsJBTdUqfi+Mzo1GaYbhWMRKv0WzDUk2cRqkFfrvz3Noo4O
mJoviwP5lxd/vaOucQOWeynjasnguF3YKdBW1zJ+WvimWM6lWyfQkFeX+5iSZeuH1u7w1+DzUUZP
zenPb5QyeYRkqUmw4pw2gXgx4785bj/BwYkic9LoDhI5p1hRGwUgYFtgA6JyRnMw7uHID2WsO2Y/
IJe6HI4VUd86zmOQ5DdHrPyxGCSTtzpZQLq+682aVL5sy52Kres0desKTWfSIUhtDEmr+TSoA8RF
KwEBOCzq+g4WGTmyLY0OcquvgbTlSL/vycuykocO1xUL4G74bAU27xenqL3l9YQxfINGThVz/8O2
BzYZ3cHvZje4ykSUWpOfCAMRi3RPrXNqDYdfiIyw/46kREXqKuIO8SGvJ0vj3DCB7Nx0+eUUYiuj
PjW9cpyowWW1ibz2q1JErOs+Os5Zy0MfMhoR/lXUpCM3stJG1uCmKvZ1NCww6Wlu7dN/Lz/DQqBA
soh8Z2Ok+xQ+H5brNBP9GJQ6Vr9xwq9UpUshcH/Oe29/OEPI9VImwGjdsvJT6Y7XO/8L1Q3vRY4c
zoINTphyJMFshyZ2o06omP5R2SX5tO5ewS/mAbqwSyny658LGmvQJLveFo5Zt+bCPum9HJb2DcEX
1byhfRf0Mj0ZyYpko+1LJJFc3yx+ovtS1n/ntNLA/ti/nGcrTiz7K3bj/h0L/489uGQoFl48Q3E/
dXWNdxRQpS66o4hUhngJZlQd7pqz1RswgFhFz4AT1htbciClrd6vmWEUQny+c6tTkXf546+MCW8i
TNYdXywlSGH4x35BOKrFoxORAxJRsGAYRabdsRSwIq2eWnhixJvf4EqIe2eEK4eYAQb0bAfGRYaP
jzsQrOWmYkO5FE/jeeBMxn9TG9kwL6FJDtIsEkJuCvZdIdqZfT2p6ytIJp2ffGzD6OfLrfF1zGtx
h8qas4f3lBoNSL8L7JaygVs49sbrhk3OYU/pLfjvMqaA7ks3OIYpAuCkZHWRJkWl4cuRYMV7ukZn
7dJsUbkcjyBMQOaiNdWpEIBZneRxzn6wrTp0fAaoHlLXZZkERh1xaxtsoLVUSR6wkiwlMqdPwhZl
ixgZ2oevhwwvoQV1LnJ9NOQo7r+Y/lwJGxN05ZD3HEfTa9g2rKjbRSTjkVulQ+OQDIH2/6akQeL3
VmKQ7F1U83MtQNlSPvchA1qOcAqzLBidPoFjhxUDn1LQQIkEqtcC3P+Me4XVmtQ6UsYbn/RjScW3
5VSJTXcwTfS6X2dIyGIkEPQ4wQEKoW7/e4PYIc80pvExSAy7wbdul5kavBzgh9ZPNqWmZcQoj+RY
IpUiIM7tPj0uqWh56lJmaK5iphqNzPQZmvw60Z5gSyikVshTYDcJbWLmUwvpKsxowKV/osdjQdYj
eziUqJEj0vNM5XUCCT12X5z2Yu9IvLJ1yQNqy/9Mmjt2ckI8GoZ+3XE4YEvelShcXlPd4mzkLah1
KkPnveKM6Np+0v9rfjA+plR49J3H1Fw43n/FyywJwORnIXxOwQ5mnlvlXYvHSYC0BCZP8jwYbESA
bKVmBfGFGhw5KOb/yCfQ+rOgPZDibb8mbaTlfap7VbMcIz0FPywABctZUXDXnDCqB8pCpA1REDXg
fo4oLTGUJj1Xyu2ybhfYDnzCBmhCdUHbrv2aSSYSLVV9V4EHnq0UM6Njj26QtYjx9RBcADGryw4n
WFBUWND4ejaIzT1tFb3x/4f2Q8wSlqcS9Q8YeBHk5haGIClQuoT/TOkraTolY1tCyzENiPnVuJg9
UrXmITnZ0ZteRDISNt/VTRsnzqMDtfqJCrkDC+xNo9+LXG7c1vZROLcC0VeJhRYtqjlMEPA1Am8s
Vgk8IbmUygHhvwD1OKtluATC5MJORjkm/Y46onwbXV5FBAcLCaaFZA25tFLY2ASbDcWRvq3ulIyi
A4/nQGgmkoYFAB4iDmHDaimgl88O6TIRPik+uA0QSvcXQ7I45r4BXIBBWfEPEmaHlgLqIT2GFBOY
uWxIDZCOH0wcMmMM6606rw6Xa4FiCkNnFfCRz3mjCD1/4URaOEaR6tcBuiz9u8jgIvjoSH3rxVsZ
CKLEjt1mm7ZzqouXp30BSPNEI9QwYF/ffoKzuUgPGZOHSEfpq+pa47Ar0lbpGRgb3G1EvBo5bluU
Asts0g0GljGbtD7M1Bd74qh+LjBwIMV64vEfaMwBeI4lRxHfWQGx9W5KTcjGXPKjzpip9qjiOViU
9Dd42/9+QzCy0m44/HNz+I0xH/9oZTpRTQoB3lkkI7ThtLiyjUPCuvMluv4M59GUVfmnVF9Wkdys
FgfIhnZB8BmXN0ZCSvXWsTFcXxwJxSGbbLGjImfYOLj9VM8Sjo6DFXUhQ3WS0CWWomij9+TU1TW+
KjY622ex0Js30HXa5hikz7+/qfl781ltsFYdQKjO1RiQUZCGkZgCyNIi6Tu7rSgEFuYGl6r9xzuP
bQ3pdCiMkhJzdmp2IOu6Wfh8xQY3CSpgjTNOzJmeXWNOgeJiXmSgAKl8uxbwn6owQeRt7SYEa0qr
jGv2A+mLxaFlNszZ15X1XXR38Gy3aWsYYY8GYKNfxwFv0D75sj6fO+Ovq2hFzEeHwcxee8fMSNEG
g1jXrvlSH5snHIdEHoX47IlFJAswbLKP/4AH+c4aP3nQ8CnCVPEX2iN3peEfAx78a8ANFqyEWxMp
JQKEbDlaRlyeLjTZ0+4LZUmOw3yKidS2d5id8Qon0i5n8vbo33bfHVOMDwAWDxxq6yt9hTbZFx+x
LpaejLXcerrGVtYmpBI1NIy2beZ0BYcURYvF1gIvRJVmkmYkG2Tuc8/MXSrVdVQz3lu2Ol9koytQ
OdOD0Eh7RToCAFieMNQlbmoYwhdA3lZCkMcDO/KLj1QeAHStZLL8AEQarlO2mwEHxWSRrUwCQ5t9
4OwLpgBBRUCr2fq4vzQQTRvNRZOYE3p7uOzEaO94p+hsifW267+BwtNUZpYVdGxhQcZoJjMZ83LH
zpLuTmgxrama+EVoeAjo3OaogWa4mMkbiv1fTzAYSPdrg16fjHs43Z8UZYJ+A90Xedvo38rm3lUE
6OYYfobL4kwFwwA/SEzE6/0a3lnflLcIdKCKWS5DJtP0BoFMUqBuwfNK8whBacuwddG4gFOK0Vkv
GxOND9Usgt7Sbgk+fWmW9VsDjNNYQ+EhYjjY/JlnNpGFio8rbpLLw14+txsW7BSNqLPFAzA3H0e/
rHxX7c3b2/H9eyDPVYGgkLh/5RFyk9njuJzxNKTtn0a7fT2ZXmDMlFOmpWfXejzcDjiMTB2B7g87
k1ebIGLgBvSC0PYihsKKJL5s5mgwrwlempVB/USDcrWuprSvKskw9ot83cy0AuM1vNwzbP61HQBZ
b3jUoPSIYqOXPSgSK3BLz47geRiefhd4as/jPubBfjqTsWhA57jMmPqSqjm92L8CZMCLVj4q1aMh
Y0divV2/7IqASLNH8OGWGb7iu6Oxr0TU/TcjBV2aEMXyJkRD45yhaWYUwewCOxFWGF40PXKKVSES
vG9kKRRzndW1x2M246fPA9Pve6wvCMGkPJGYRNQZsZzenCzaNhDfM9Z53lSl7QLoAtfmQvnbZuLe
6n+8JmX5R4osR2dQSJOmyHOImHiH10RQtrP3mqy/jm1FSyxCIKIcieFu0+DAqDP3SYd7ZI36+EQI
AvNSt7mH5EbHTXuQwrWPVHiI1DiZio0/TvNw3fiOK60jhexsJYZ3Bak1rsdl38nUTNeP4KZgevSG
3Utpg1hI1nG0oIHU9UpSNDMIP/3efS/uLdppcSK4sZ7TmIp8HIg7oSdCEVuUis8H6WsNgkYyzuR7
9nOROeWHtquYxcO0Uu1taXcBTK+RY8anzNhVmtLznjoT+OGCjEZz/sI4cxdZ6baBfzXTxj66q+RL
diFCo1vXyBMqkxf2hLyI8h++g0iKKg9rlH7ZMT3oeuD5mLxxa2dXIrhgAFh2TPZL1VDetfAvlnzr
o180fq3hbRx7JIIgC1DwfQYmJ74/6o1xcwHFgk1v++y08JqCjM8/yWPD5FDrWUio7i41Cbje2S0S
ZVvWHcCTo+Wsb1fK7fBrdLTxr5YVpdoyrTn0lW+LkbjFy6AVpiNNBcKHj7XlW6Z6hpdic8IPR2Lf
R7xnEo0L8JUwszi9ACbQApXk6QRok6rA+kHb24CvgL+lcRQRolP6yJOoBqzJEyabfaIF9hcYOgfe
9ek96robT9Tp6RwTsweiW9usqGJx63mM6CETJ3ljFZLyTNV4yOYPQrUU17QCW8O8W3/+QVR9MAPj
VfhVdUUirnkKaCo/QBpb7IloANl60PHN7HTZmC054SY54Dx28EtosvdI6yzwOqSbbqApW4kpT/yy
+H/l78u9rWDd2iI+NO7YDx5bEEJEbymnifeEQiZidQ00TI0j8y2/uX8KKgvSQWvo6HSstdYY6hrl
mZQmHlchNpoOamiFNo7kj3QlFtlytUP2UbgedevMYLfrdY0T1vSqUlZhl6tm84yuzYNMVU4bpTyv
BRieh+lYEpOvOkzHDW7hSHISf7kSYzvnXuWZ9YvTWbaCYuquCTko9f5W7aPU9BqcXu7Ph78bYUw1
KzWSfG6E/B2fKvv/DRR3/Acnkygtj4YSU+FCxlXtylz4EudGSOt98MKehUDEboUTg1Hgd+sfNHQi
07Mf6ActVxjAmMOORCPQ0F+bkQkhYDzM5jF1m/jmSlky0Xehl45ZUqPuY47Kg8Otpo9VS80bTVHp
uIFWXNnn2XTRcrEbtAwPTljT2diq/0+HrbbavHnLV3g2CPJYy4X5akfU22myrASqKB9Mi9a1XbVI
iu9eXLnqQhT8ns1XZtTLdJ38zuW8u2mlOs3zdu9si8W5VsiAu3EPn28h3Ncbbikjepppoj4rJQfl
tre07YizJQaTKJKTw5j3CAZtvQoPBOU79SEWDzeDS9sGMbrYDZfzzKyjpIkP5j7Eqa8kNZ9sveT/
YT5cigvIehaNq0tPC4DEgu9VjoNWUtOmvMCVXA3UfUup7IHSUEJlYSIHfD46FlpvnAUFOhAw5FJ6
DauoVjrm22VB2pweYjMGSJlNwed9hYTZRKzKKzgjQGFNTk2fUAUuh2O53G4iToflqRQERSpd+lWz
OctqdRX5vvSWMPp3gye7NNWrpw6pBnX2C+Qd0kjlSBU28fa/AwfH4j2EEGI0Kf07oA5YOajGI0Y+
t/JnxjP/to0oi5fnZ1Vi/od8cCiOi2uV1yd0uuMWBnmu5yBaaNJOjl0Hi/sf9HK64XPky2klzMFD
9MWcD4oHPk19TwHbxpGC9mdEZKPEJd18XX0VkXFnEE7Svf2r01g1oHiwgV1VvUNAVHxyh+Hp99lO
7Dfd8mHQP9AuW+OnkMsBx2mN95brRb4PSxz3PLv60+JaU3Od0wwMFekMnkKw6zu4kQiu4P5QFym+
dv1FJzu2rLd52Y3CCWtK7F/vMXwjVUujzcEGDBia/Vs7wxjmxofBZon1/3Irnki7ge9miWxElLr/
3OFe1kwj1gRwG7zwzxHH7bfUOLuxFRm/IvRNBqQIswrR09DrSpwA2LDLDyDmHkCTsNK5R3xJRn+U
9IF61HSasMFh1CtjAjrl80zWJjENIuXVARywd9yKIOrzeM3jstXnnKbchHi3mPXWmK02OFK9cJdp
bep3N959Kzaa5BHyguoh0rzyPtSPsOgUyaTlIhGZFQLsx4WP9QKTEZrtwW3NQszPcECGlclz1FVc
dsX8Zwcwc8zSVL/jPuMmmdWcbpJ/vRUf8s6FtbpIWdwv4jHBzDmIYjHPOZwVZr7Ysn7gfYduJEQM
y7t/1UYttvRtaz5kyZkIoTkAnvWsbb2iLvBys2qG8AKbfhhIV4Q/k7ro5Ie313olC0JoYeShPcC0
Um1ILRaL7xM7Ocx66tOgj9cMehuHxR/KdduG/CDPrrrAcDFeOyO74sQIZ01c5PpHDaDQWazwrDEg
3V2j8AcrWNIsEMLgLwUm/6+CF8cee1AbAnJ07urOw9GVelAoLIiMjE6fCnoBvUqvCvspZChn43to
GPGx1UE+xYy7i9KLGWdWshHiBqIwx+0JLDnP9Zjrc9XPdmdbxJZnmRHYSk8bsduxgKJLWao4qQGy
D4vOXr3XHXm8k1BFXzl8ef0BdWTPcCz+LsP06PEPBIWp4/qXMoSNabTxfNyRMVe1vcbLOveyuCiH
bNulq5j0COlWqowX8X+SjGOtqkWTv4ecgrqXTyb+g8UcISAwRxO3SpCklGbGrLMwUv0yMgfFaHyQ
JcFBxldsySZh9ZcsDlo85vZnuv3kF4Df3NLWBQf1pDqsHHgkC1Rh2zMPtRvDA2DceCEsYpKGNQcy
FDkXOsRoztSeUXJji7NPrcq1uZWw8/+kjUbKM8LO9LWcz+b65kNqU+GRKUkNn8I1Dsxh4UM8mBu0
lMpdhECdHBZ/Pi0wYDg3CW+6iNG+dj7EWLfx6uAaRJfciy+Y+GFo3tAxP5Pokw405PHeh2jnRxPi
7iLK4cMvHRm1+dac5Jbee5yLwZUNkI+M/eAttu7QdSK9wwUPRzFnhpDyCPIS4JVLa6ht7U/SxqMR
apvQ2yRM0zq58hP6YlX5Wommra6/MufgbmknbUML0zwO3kKvA+wJFjJiwoyHbueC/Iz3N2vcIQ5j
2bB8BHFI4miK+f/eTr2d5pRdfbA5gCFXCGLnPzsXXFZP1/lT3Rp8jIv6Ah5fDXyNKIo2Xv5tUcUr
UYcj+gZuQllor4jQX2H9s9GRp4/yan57YkkPTMfHYxC39JQdQ9M+b21PqHBX0biDf6jAOXMPHnqs
lOA8lwfZMYzMAIzd4Db1Q1hCP0q7N587XgS9FKVcCtysVmPFMquLXCebXpxN35wIdLcYTNFwszRG
vIyyoCxoyaN/Er6ubJFYwno0Ekwryu7xapYi73khRVDdfaHEUZVoFoAgzhml1W/jGPcsMMZIUdr0
HvoB5vxjAn4UqbrCJtohaWsi+jo/dXkN+9WonfHNKPz0p7ilKiG8Nu95jmU9UsYSwBQCctmL2gIS
KFzcBhOa052C4Mp4NcwqtxQ6YLbBhDnT2+obOSviY5x4mfWlWGklRKwrAZ5i/3GgITdy3Wisfdr7
4CcFzhEtxNmWKdf+P+DR5zQRJ5fqXOOBIBpYgEvSRgOw9TWX48OJ8FANyIozuGjxQbdKyCdD3XWN
aDE5o5oc+Ipc2lQ7x2BYA7pQdodPNDrrr8ZcAGz9FlQUGrMQQEKKkaZ5WfbM0cOIlX+EF9xtgMqr
Qj3K/+TM6KAl+hXIFDsNQDkFEhisIrQQQ44WMovkAVBbsY960GPTXU/pAK+mes22AccR98NDd3uX
EMoh5gPRGF7qY6w5up6cPYiGHo/r6dNBJOQf0MaD+gFW6kOqnO9nZAixfZClP0m8wuNyQKYvYv2z
WXrX1kUS6JAHbIAIaRM/KY3Jlj0BaKodGjQuI5frY+EVFlj6PtXVNQBQZMop17zYRweN5dzoFWfx
L1erIUxpGWUbUoWq+wJEhhl5Qu6f42QSsb8CrFD/DwpGLup8b85lKOMjETlVO3PXLiJQkehHPA9Q
3Eep3lok7hLSOPknkx08j150qqxCQVsRC7OmCKgWOXMYi56E7h9pCOrK9F9kANXpQ0QmmVyeFXZg
i+W7TFwTs/PnQCLFwSEcnMOeLCODsa6odhno+vjhJnWcqBUEVpNpmJHNKVHaIM91k9fSdwX09f9b
0P8xDf8asnBMAy0coJmqZ5LkDhjoKHuChdSReVBU60lDa4pwR9Kfh8e7EFq9PCRGp49KIP4jy7LH
qcCmuOBmRDWOCVWmlBd3oPaKgB6mtsT3tLmYwI1fRddkdBM3DXLLH4SEVt4kpEIyUdWzyP7rPhXo
hpFjSS1nth6zFA8t991hNOV8f0Bmy2JJZ4Ha0IhhbioVDxLTjf3mEa5h+MfQH8f7bMtzP78obFCZ
s/cFqgGI+1NpdwqUOV0aZLexWiYhlC774qN6Yi5oIEG7Y/VTLDVqVvmthRzelabbSeEpdB1psRyh
/v7YFYNned9vwVs0K/BvGYdJobyl/dxBzYUgjg5D7MvcvjxuZQIFlqV9DrvWAo3a7SQ/D3erkBvR
KQXE7ogLyWKyZ7Kios6vcXyR6qi7P4jhe1pITAX1ySHf0EAgNCn278mfz7zQ4wDhxasoXeTMkWyO
32YHX7BLdygYyixLC288i/4M6rm9oD9a4bsi5QJegHgt++yDGS4SGeB40X8Z2VrdlTVirU8iqbw0
aqq9LHDhJ4LDGfmYQ68gFLrUSfZYEfoPxGgIZN8cyJvxgsfTzYZCcOR9l3BUNME0QUTSCGEgAMZT
x5yCsK0OPD8zBskWPdnjyUG3nEOHqhi5uxooRT2hgyn+0gCqRrF4okp0LkPmyiI3KTQ0iK/3VSm2
JcGeM/n6hGZ5IUnLxDrzzoV9kqiMJRng5ug9M5Ta7WudJZuz+EmiigY8PcTkipzORpcB8IMI0Dq6
8mSBQs6Xehc3AVNmdDq3pVnnAc2SLcvYEfbKE46iTzi3/6ixka8ICd2BAYHzzPQvHgCIJ484IEQV
Fhe6zAZ1QlIYEA98KQllfEW0z3AtziIpqJvK1FONRvI0g/++uiWWk2yAjBMz1sraA1cSnWshPFFF
6+ErVbHZUqJet1bMeIcaeKrx5qGNiU+MWf3ewBHJoRWziwohPxQJN8MjU+MbAqyY9CiFek/g0g/d
yQzHNhoGkBFhKCj8LBXDw8RDTQNYy+ldseKlpvtCi29xVlOfFbBANnclL2lu1d9sZXEr0ZHUHTrw
272pgUPdsW35CNqW2tGnt1Mf+/SUVFVGMihxd+h54D+z1HOKzn23b48jA8nAh9gp1KA3gj7/Uf2p
5HCvNb6dwMjA9ieCuDhFJ5dHlshiox2TWtXuLLSvKHUtao6OV7WvubojBDVaSq+bK+OtEgvqqDpe
0M6zCzfz4BG0CRhGwKgNYmlP/k0TneZy47FlyxxO9QmO4klTdtChxpPkAIj5VWnG0NahmRO8PHHI
0zpXsu+f9DKpkOmkqXevY4Z7wv4iTpwXpcRvJ7RrM1WyzD9n7ApXRynFZI6woAQwDs5jbd+wxvJ/
JOmSqD9QECapOsOS++HimJ6iJgPArUcNHLyLAtARa3Eko6riXQ/YSvmU1cIRVoECuTqbxXNgtSvR
dqfcvGdgLV7WxgspD46V2H2rKWFoA18nFZwSm7//kfi6sKTANRHH/i/1stDo07UDuX5A2e/aig1c
i0fdZ9pqTZevWcmX1ttcdqWUnFAHKDQ16rdBCO3Pb6tJy3Rvq6LiT20Lzp61Pv9xzUNjv2PQJF75
BbvWH9tEVGJDfwKkqHyKAv2lV0Hj5wcWyh+MEUtW5GTVWg6iCWydcphgfK4ilU0GYouCvCxIz2jv
HQVpH9LuW9ooz4iDK+LtBBfWIlI46AD+qMAh7pO6UPa3z78ztjCUGB4MD477ufcnLURQDV03iZEL
/B5IfLFsGsKKT20SxqtzucdS8a0Uy1VqDO5idakPD2PGBEA45RiH7ugz6cEguV2vUqz0R+sGu0AS
euMXL/vriUt5VJ2N1XJHkYr5dpL72GLUj09pYKSKpHm3z+BBDSGWRlX5uAw3lq131ulSjZt7pCyn
lJ4+1V7P7f2v4GOYhv6iLlWGl7aaMxd3yYsIDwB/F/uy+nQuzuxoBSK4rVnxzhBB7BWqmVt5g6Td
Ys/334aMgUF+7af1neVF0f1MFbEIJwjDgzQCAw59QFPuz40C2Ep08Cz37vFtFYPv1jfLcxXfABG2
7Ztx4A/qbzzgM7zx7uxmrEXp+IivElQLIZEEcPhYZe7l1zurkKjY5cZpMDGgBnewiw1WQcFjyoOL
BpkzoK8DEv+iWFcKBzOvOdmgBoH4LKoTM8TFsVGGHAN3UCLfj1uw7Y49rmHYGT8bI+l9lAY1/M7b
yePYLOP5j0MFceEsRJ1rYVVaDPE40zIiMAyJQpXbQoB1aONT1CsjDqswKmL/YWbKe+Z7rQDuy0Ah
LfO2I7FOhQHMqWUqKUCxGSmHIpFAjMIq7J/Q8422SrooWN9fuvtzsbK0Ls/KowLjQc0dqxNO1ccG
35swfKzBQMmWcRMKeq1N5lF3KCpQ0ZSfduXoMPtLHvPzKGACQ0E7iMZKF2g+chOiZfNn+A3dTIIC
h/50sSZu5MHNqGU49LKwIdkuOX00jBMTEZLqRA9eFFiUrnFLuwEj2027cOrUXsf1RugyLLfbmnSY
nF214UR1l1DZ6zzoMR3aIfqD8yBHkPBRixDa1Herru4K2IaXolC1vZ9uOc5e7l5+JBnRRLzY4z1i
9JE0AGqPbeGeduJa8uqrnUzXTsDzG8T/XHCyqWEzDAxaPyzOlkBH6+25qfTfkjS5UZH46ePtWd2j
W17yCTUBDdP1omazCWA75i0p5F4b17xqh3FJyutLm+4Si4NTE/W2WyVAxpqsKvfQE+VPr+ScbOoM
+Jgo6orZT5299wFt3Fu4v/Zqa5oCqLnRgAfZaVKHngAsVx8Iq91uKkmzVoI+8BEm3qpHOySbe1Lp
US2FM8xNzG0JdXYruSeSdLKA7lqTnQ4CtaGpff89u08R4nfY4WpO4jO9Onq2JulVMttvIMSMQvKQ
qlF1pZP1aw2bqpbdmtyo4+KSrhTpepsRU3xqaJVjQB99J4NyThmKT1qeTV2JCXB0JhocgBAP/Nay
2AS00ToMCDSqheOauLPW0MzSLwB2zS018w10UkoGjPAgnvzL4PLSlfqBNkrr8dd+5FyIZriMqSeY
KdtTPW0e3D3/qPJbj1JF6tFOYg7iOUOO0vmcxrddzEWrRvZVh0hifWHrNQcxhaUVP6HK6LUVfyYL
SCaLgNMbjwmuyZQBfjxcAIvnvyr4eHgWx2a9pQBiZbmV7H3sx4dEGEz6ue1gMYEyqRNBk5C8ypHY
I01Qk2Ta/jkdzAEA/V7gsZr2j/5G7TkQfwJGp3uCwD7VfjlNvQWd2apd2DNq+ixtuzzr/o9LWyZB
nLy5Tk2W6lcT+njaLk211hD1BZ1qHViQyzbss9c2/MStYlkZ43zFeNqQaZTZyzCE3xY4oEtgdJWg
y9OA1yvkEe6NNVPgux8MU2YskAMyBO6Gk89WoMaObTvy8mtA0/W0GDJ/O03FLLQ7K7AMDGghF4wm
7X094ZGwzLgM5Kzc3jQCmXjUM/FwNJhGSbDy0YUarIu2a2z9o+mxzsnLTnd36CC+nCcfpYK46ppJ
fbNGrPwdEyyJb6Y55kf/fmfGSy5N1ny5EamFb8TchHyE2TO3KeW9Am8IDH60x2LyiAiEfrvdHui9
Ts4SMCEw6zy1wS7YRUJLkveY1/31yG0UbyKj5ZfHDt5tzXB4gspBxeOQnSXMftdMGfPdG6vRtjSw
PSfNTjuaDTAMNUYSWYMkq3y2UWQXQSXGPxTkRJr0YqcWR+s5UoBQFttKYS1mYc92Ug889ott6jNr
+dgTBh58cOGmbe3qSxz2ATOxx/x7bRiDrSMLDntieAj8TvdccCVIIqw+9DvYuAESxPQFbtpIH8Na
2li2JLRTelvX5YaoLAqczaEgO3SuL0O9sTWWTczL3lf1h7Yf+8b1F8o8sJzJEyEIDcw9KAvjyDcI
EZc6de0mUcnYg8CXJ2lrN+YLtKCABYJSY/ZXoKajZ4iFwlHHLfGpRDHGiILaCaEEylHwLQAvg289
85ntju4c+SWhp3c20ab/cuNwEXixvTCI4/X7/tYhOAkBE9OdeL09UC+XruM4OYTyuiLyYiWySE/G
fPsBfdoSeb8tKiNBbx73+oiYNDxH6b0mMXV0xGvhSS8gNuqw9hn1zTNKy1Cm7hsDJU/hIuS8Ta8b
3yXpX/bey4wabFP5Y0AGrSe/VYsnMLwYf1HRfdaW1xElgjsL7+jjHWUiO8EfzKkBOg6dBlvrsbO6
164q1TYbaFOuX7LQDqSnhgnlbK3HHZHmaJJ/yfZFQvwZK74DaX7vPJN4jdBqj1M2WXIuDY8oXfot
hBL4Fuv+XJ8kawVZuif17bDXBGPsAIQ/8EeS2Xx39qTyELfpBDVB+cAI2vvMxNvwA3VtDD6LQ0GB
9G79Nn+enRM5qb/NNsZSAD6Zn4CfIcbcNcjv8ewv5QDyU9OjLn0rjSCL9ToafUYVzEnhS5SgkajH
bkpPmtkMB68oecJQ3NpgHbQ+XZZA6xL+Xf6Txg7/pKijYAEo1RTViPHeRWDpgComU+h8/eNP+0kj
6I87nWdCTl1KtkRJYRBhW9JP1qU7SX66d9I/DdLvNb8AgYJi3b7y39Nup5TwXXprVNNzBcViCoD7
SQj6LeDt18XcsKlJvh6T4F9+pC1okOHUVF/PmdICsSEkM9WEWf4Zq/vfAcTrWrLoraDAz+2Bz+dV
R7siG5XTLEJAcF/wHJtEywA+DnehLGXj5Sry5JpIP9Lr9xJqUR1bmzAhzZOkDLet4de2lUrctCvF
mZIh24f9f4ukh1ZIvyOHQ01VqUgrpOAxjSXFTVFXgY20UhhE9Fh9kOjisQF9pn1GaawFhEldmNXf
KBgfn5svSQCWqeRuU6yoHpnLhwf8anWB48zF3/BB8hqF2AX9TTnwq3SJ/L77VzeTJ0Grq3s1ewYd
BGQa5FmgQ0Jr6irQzVTJXbXxvWsuEU4yIZSie4N3S7b/yReFsk8ydrWEVMTfPM0WNavwX8yM6f3J
ZoSYwPN63dbRfJ64bECY1oGob0+GDhi1gdkgIVlRrAAyOhJzHsAmcPnV/E/6HQX38OLJqJkjpRwo
fRxUqjRXzwOb5KhPbLhmBnssGl5jp01/zVxJIqbWwb+9wSU+iFCkFZ96WhQNHqjJ+XbHd449wO/d
xMLRU8Fq2vQBxb2/R33/AgUXWthVEQkVA1Oueg0KOvyFc82TL7VWjyhOEd9k8FHu2SkJxjCUGmLh
/iXWFKSA3qld0PSGCiDJFC1SLsTePm8AIX1sacGAk2g9kXuP1uKQiRm9pewqShwBJsTSK2U8NRSu
OVArEYwsF2r81eC9vQfM9+eA0NhlwfvaECX7FcR+tbR9deWiEmHMN+P7XrDS9GLVBDQwEv4EeiaX
gm47GecI1/6qzjOXaA0M1dWZkZHuduAduSCTZsVEaKaHRghIi3zLNoyClj+Xn/vWShQezFXrk+Ij
FU+labIeTwvMfENTId4huR/FXivkOS8H8kOdATZRvaB1Aqba6gYabUqRVfyXbJjTiozp9g/Cm7+v
H0iYI+CGoXkycxCKY84nb1csCV62NDze1eZxgUC1LiZFi0nLVqgyMAcQrlOlodoOYZr+M/MePfuY
p0OJa6eC4SF2ncEkvIzbMGz+YcxntAYTIw7VwetpUuneguzgTWfSXZ/2w4GmIffhlDCJd5oowDnn
8VLIS+kfyZufr1bgkTIEZD/CPCXdeyaeHXWw+P7PSmpOvAQgw4XRJGioQPod2dTTC6U61KFpkl5B
xaukqBM0kPNQa7IcD2DkqyT/R2aK64g5OgKCVjcgmavjg3UayP1PILMME/GRWD91fqfc+dxWiSYh
TjjI/2Rr15jGAFRa1sjGASlLMzoBTad5rMpymEwvwHvyHZ/M1L2c/pvwStCMzw79nydi/YeAo0HF
kAC8D/uqvZTL1jpwXaKKNrUXzhV2L8gmwD8resj1gA2qRV3JxImZXyTe6ZMMptIgIV0jI1ncupCQ
WH37cXWG4dCRa1takkgAlvdH6ChNCoQwVuZyVYOs8GRCyu4T1+atTtdC6V9/Hf3BhrDROJpBCHoM
bEKSXOmtvKRiEEWaKgoxFUfg2rZEv5JB9nlyYsTzl9ks6ALbxB2OLT4teUjx1w36lYenrjuOMyDj
Y0YEajrXHcQzX8qnn9MqiXpfsNQJEnHmgVoo0h0iQ0XpqLPFAvAlD3bmnDtS2LTAjobYk93anI39
v7kFr5Pe39rWIXm06ULaO6kbcLzHug2gHpy3bJGPlx1yF5zcwXx3ltvmFBX9rLw5G/KvhLUY5N0R
h15EGFm4N1G5B2hQt7PdU5onTdqkU2aD+o99rKh+L7a/8Gsp1NRXBinjt0zmRToGkowm9Y16dUEh
bcgzqa5OCjaO/FCh8Uez4NhHsWR9hVlAqjHaNkeJLSW4+/nDybr5ypUPXHMRBw99XHIyhJxU4hLf
rD4iAQp9VP5vXC2ISSE7qtmGFl13cIvs4RUeASNjIb/EfZa4Pl2sU0W4KfRFbk3CMupw8Chn0Ceb
35tWMGr75c2tiOgvHeosKLKka2OLjMMOwEthMy/QnS8SGcmXIeFlvsgDk2GZT/rycZ+71S2jDiac
dxvxZPxFlriLHgJ8dxxlTiOqjXQ5cCyVweQdw6kYt1MTint3An4grdmHK1BB4JihdNaObntlMWFG
pGIl5PtVWADZOAV5iJ8GTUM2NFa5gEJiElNS3szOE7RAgMjXrI+rsQkq1ZPYa2XfFr+vRn7xYNgq
ZVw6BOvu4yiiDrHpKo39vdAZj7hddHxvMzMAefl+R9xW5ErQh/SO+Fi1tyPy2sH4n+qMdJ70siL+
vloyczw6RiH9UFHZ6Y4iTS8XBoy55YTdZ6Cpl49spbt1+R/561spzSqJ0B/+vAplGK1+IA9Zwynm
rSEQIfaDve1mPv9dq2b1LgIMLsoGrS+/laaxBDUNnRlpUmwLoFb8Q9qANiwh9N7naNlGco12L5vd
HePe603r++w+Vp7SLWzhlJl5t0Jlv+IgRgmv9KYzbYhu4qlQAWIGTXkCKbguUPyFCA3pWWogKpKh
ia+J4ANRmNRksR1FGh0zX3mzfZOgotuaLHGVBRUp9laGE8mjDQBD3m218WKo/tP3S9YK2+PrGbLx
/GCFyPIGyG75Bynqa+eeJrfx+1Gbk4ZaKKsniv4xNceBz4wLZRexpasyjgozbezEwjbfSSHhPVun
vh3uRmmEZxrLzoiOQQQds0jEDLxyu9u9OlpKpBXlkqJmTQC9t1Kjh423/FLITeDXnOwlhfA8HNRp
mLxQsv3Y5pk8r4AKfDM0uLVIOOxWLSCGa8hSRcZXB9UAUujRXF/6whTnSFv9atk4+Rxbrmmvkz4w
4mN97FOCXEDGa5kXn65+J6M6bR+/LDDAKiyOPrVke1j2KajDY/rjUPyxeKKr62eeOIuYKXBkIpvL
Yv/Rhf1qkud6in+QR5boToB9MszJV60iI2dcgSDvvasaw355DzFVF9Q/sEA9tOL7JQnlWZ7qY/O0
BOjnckkBIN/WBnEoUSWMfDGNTI+QVDnn8U7sFf8kEbN5S/BDP6PYJJ2B+sw31EPEEym4EH9vrgQr
mezMWik8nalzrDcua4qJtuuL9IlyGvA1qIOs54U82WkpWKUB6ngysraUeZOwGMnjCrPyMYf/SIDS
HQIRpjqbuh6lMZDWzoHlkK5p7Cvr1LS4uoLs6dDVNk2692Nr+GnZmKKCxUG95lqpcM+sjTrM6NqI
ZuH4UbbIok1SgZY5h1GhmEHAYHCKCgx13fp0XumAxvlQZpATgKPYgGVHiAcwzjhRIrB1VYEeARj+
VenfLoKI4nBg7hV2zeto2Z7dsGICphZw0CNOfBU7ABfy7FnRs5TSkovnhuyhcUGkmGuLEliaWo0F
PdDLymcOyQ6Gw/krdLQx9udKswGXWiXeGO39z25rD60Bl9tN/YtTNdKqJtb6aw7JAihcOdWxT0PN
Re1O7wEDuAyOpCSDIR3MGyEVNhahA18tzPXuBG/dajWnTrRiK6myjAzsQ9DbYXia6KqmsyHQEp00
xJO5GJvxNLrSl224gOo+LeROillcS1FQhstdhjso7bimzh4OyspUpNEbxgrEgRQdOKOnh+IenFsy
tXcqpfocVNAM+vinfzGtzR+0GMfnALXw6YRgR0GkooOSMk8pemKr59ytIe05z0kiFVW6bMS7JvNZ
u5wtdWJEQEb5nvNj+vfB0wN8pXs0JyFwprGQoFvD+1+WnzAhsSsxR5cTlqEzv7yyN2eKUeP968+A
86VjpYBtqkmuA5PIpqrFxixdTHI0hqx3PQdahhDyokUZBtI529Xz13V6EncLFE/j5w4zlMxg7tSp
aNQBtUYut3UqleOzETO6o7w2MOnbHkVrbudg/z0abvWI8mSrsmbUqaDUeg+FoWNoYQvNIy1SU8Y3
3or+oK60DA/axBI1GRwSeLE9hm5XUmKD5u8Tue3Bb46v3n6VAIXCHDKx2d7dKqDiZRWrWDBJFg6Q
ZpmkenC51c/JExO0NHPTy+2tG+IFGqfw/QoVwT3Df894toUFxHSv3FTU6Iw/BQVZ8kgtan1FTxkf
fNh0DFa5KSrHDzNP4HSa8cLuVief8UgmMB934An7mlxZcYstqpNzvN1/etccE4YwDP0eBB/pQcqM
mtkbYAQzrFSZNEsKJ6ByMxX7kRAqnMlSYiVxpsyxYB7ePsz0X6s/7iTF44HCXxQMh9k3sGPfQqDB
FYxO8B+J5Tt75c/QEE5j3p8tg6TqHciJtLWAEcMZoOBK7zXpM4Nun6DAaxAzaa18vFDLxj0YVeDz
KtFa5doM/YpwVm/XABJxxqUE3PyHScjZcV2rOKbb+fw1bOW/JNPoporuSk4FRQtKCIpQbSkPf5h8
Ud88JMM9LYvcJVMb8U740zNqHL8+zxDq7+ujz/CQUWFOcoUKEy3W8L/0IPs+7oqTUaFCzPYS0sra
9UViytWQUkkCaJrh6pi+1grcd7fyZUNrldz1u7ACchBvARRSXCBZhpq6T/6BGN5Lk3lxIXgma1wU
Wm3zFmYkIqCUBCAVpRpq7d9O50psuJ2kcQD9K+ao2WUt1rrZyqi8YQS4D/qH+OAjHsT+6pu3QZTe
0Y4rJ0q1nRwJfYYDQ3kgzXqtZifpcJLKrhokReHlq95XDAYWnXM4HHXtnndlOLAx61r+Yuz/APHE
ZKSLCwgsCe/Jwr5xCrmzwNCnigihM6uoWoL/o5TXcPpu9qNX4FuD8HlFg0BfbN0l4c5YIslr0BcX
MBLXDT6KudqDIzUDl4psXycVpQGzqkos4VscS3KAgMQ71SAl0GsJGyY2ak5WGW4zBfRklwkZ8NFC
8lSU1aZ7YAGzZgEKPQgSaIPflS1JryrX5KI+QCGSDJtw2d1980DMvHnQ/zyIMyK37vxyMnsQ0LHv
h5Uvt1WGjGByVWeh0gj8r2nYxNZjH6IJ7aNnvL3UcT591ANqIdczlWdV/uaP1ySDHJGDkUMg02G5
7AdruWK/ucID2zgc3oHzWSioEKEEMOwh9BSAj+ZktxPCDAFKCiizbVuhOVzytSOLgDgHpEOCTHWq
iM4L4ffITOdlNJJp+qu9gP93krvSeejw5zRLEMVpbITxcnnCclU1BGoJ4Zw0MiAWLOQbMYgDtM14
Deju152e+cP5tKJ3PH5X146yUklpZqS6K3lDLIxg8gs5rnjdDTZn557c4BSfN/SsHnRmj1IiIvNy
eEmpiYNqfMc7aFiS+vDjgqSkJhP4khint3JNI/AxsLuPu0vscUVM6JWUgGwFD8PVd8CD/UEHMLg9
vbPRmeBlJ//htyyRsNgPdqm7a2gdV6IM7UYjgaeyfajWAZ0f+ngv4itLWDi/0fplCZBdLEvo1Zsg
3C1x49YxCnJIvKVXoX4aw0C+Um87jmQGlXCCeieqauar2uwaiEfk5uFLYJDO931+09HXOj1LXKt3
Aq0rb7l5H4C0x3CKjBUKnbMJ/UCYvdwTUxLd8erYKiIBAp2X+daFzzTY99Y15+KsXxiiMPtQj0kt
qH21FK3dJlyId+qNkRhoO9zMUOMZShrnomei5fT8pANZDfPzhmrnv+GHzTjEXf1FAHvUKTqFUUh/
FolJH6qwtZnXvEAKSBJ5ZkyEI7QIPFwQI63f6h4fhzCdKaCAKG6n09Oq/rAEbBSWFoUVlD0qaR+S
nZBdH7C2Jpz+8A6cwOLfXwZ6CMP5ZdqVNUf5cOBk2BwmOnbk1HVPTDB57bvWqxPjb7a/JmPVNhtw
f7dILavDVkELGiyWcPyOY8H4Yo6Qc86w12j8VB22LACrvyKfccJTDe4mGsvkdDN0PrMeaD60ss6p
sKTPWNqGp/UQhM+7kXmM+/mNH9ORmWhU7SEvQKUz8qGF64NvupMnPl8V1ljahXnoE01neG9EqHby
8DbGLqZJbNQBkpzwW6QktDGsTJ8Be2CzMFRiZ5GmttMSVaZ8Xqvb1G4gca/IllRcXpV1FNjzNCum
zCVKS8In6jpkymwNzoUKtDYnXtV2kZPiP4IRi3SxmbWGiw+TAO4kgt9g155Y3nNPekUkKHu0M5fh
sQu44RbIgtQyQXn2PCTgCdnoBAknLHbpiQ/5frzJTNtqxWFTUplOv8fWPGU2ZKbAwtCxIKZBbOPx
e60wzcElVlowpwx0jiR7qj+hcBKBbyj1OvNclbaoP5PwJ9IkgzbxOdZQaB6nXEZdcdE6/MxoPmRP
tvlNMoUo7IyaTRRNY0pTMkw4RL6gw3pSN0SAETTFe4Gc8BegpQKRYngMUkXuERshFaiKrlyGteCQ
1TCvS29pcyl7u9kkm/LkOFf9QKutSgPbiSHGLlJrwWYEp64DzX+zdztdsTNNNb3Rz9ONHGg72kfA
BUamHrmEeUE3NhHMoe8rDxb/nGrk7Xp24AERW1v+2WGTFylNW+CJqrLQaFXtykcdjmYSoTcsOpUv
YozO04Yu3JAYz5MBlc4mjtR4Y5FVWjCxVyDBJsDQMomre4CgGA9gvZ5eYCCJQMBCcl1DTUhFNNZF
eoWtUAjucG29PmsWcvD7rUK440jxIDUPQY2GqYqQGuKeT9o9xC6Squm4i7ZizjjrE0rQlGk3YQth
MwXRnrNvzw6NXkCeTRSTVqE+dsMni85TX7FVmnjg2rSTyYtudCczlnsn0z+JmI3ri2CjsLKKCOZA
6ZpAkUsIO27BMSvosui7tNz4DiEmmoX+HyvFx+zSjX4vzlhf7dYG6VXm1Coug8tuzdIDXVghQ52l
gciPAZdTsM/c1RWTkFkceUFP57W4KrQWCtaJ6VwyEiMOj6Hfq2D5PLzVHADoIu8cUecL4MiwyNed
4vL/ZycFL16NN8cw827kjzT+KHWfkqyxxvMywVF5tC3Ax4Ljb3T2yfYFGU9aF6ayQg9xUw37CBnS
AqTwTxXKl7Uyy9QUIQaZiXwjlT0Jx4Oh8oxKGkLu3uO3j2Gdq92IFs+qxWdwa8ocKrhlWK8qLtMf
K7diz3j8rsO/jgWUGDAVn1IiArL3dO6n/NPfgvkOMmrDWCwktfeWdmKPWbSxkzqP3XeY3DiLhsHG
2ivv09nSeQLiixbWCGtLI74yGM2jSWjd4MzlmhEjB8rCe60uWyUo1sAzfsziT6bP8lYLASYl32Lb
WC7MH2EAFbsSLskkRqK7yxrrJmx4lF8tMn8aBciqv8gD0lXADNkbOIjyl2IEyl/R1GSRIP8S2rPr
9I7Hlo23YMvxrd1eH/BsjXvL46QYC0P0+nVjRLIjs67OzRSmwJNKK5W//3+xC+lMKccVyKClALdS
j745Venc4zSBBjbDMrmxw0xnKOARbKXz6ZP8FVyh4/2AT83C016R0PYcdqoQkHk0nb1ZqfEcJp8l
rIGfoSrCbBjNf+r8nWwmL7tuElgV5gixwmcSZBoS6MZMcq9FNp2k/Ya/2hOGKwhd68OrZgmde5+5
nqZYIg66YlKIUE+xanl+m6XV/Pfews+V/eCfvWaWR3+VfjWNgDk94xRz+H0v3kyBpA3pOlmhECt0
dj2gtuNnguWdaGHTxvzZt7knMfW7W+BAUmqKGlN9s5uiRFmPkoTS04QBbdAhsGsYMzUgVIo12DU9
vXTZLRr5R0uPY7PpkqDsARouZ17F9tOabvu9Ayd6bpk5Q2XDgO5c+HDGUZX13CuSd3dbA/y5pnuM
I9qRjGawAy3Y9j0CSj6+UYQWhITXAp4YTRgH5O1p0Tr5KE+TQB5CP13y8ujjac2FbKTnLLMHca1v
K0Lq7fFDKC2IurtSs9Tvsjlu7nzcBL31eiH6n/KbRsgUOvb8De3/cvZclRfZ8EXMB0q8CWF4corR
jINXu67rH2AglWUg2e4LkSCBQF+23r1dFrJZ8TKRsjbaUudN7ITHF2xzs/upZQ3Ls2/z7QsaFTlx
MQI3rqj0sWoHoA04NsPcPduRiu3RacWUsPpwhRSxag0Q/t14wUtT1ogrgPCuvpNgmZtNjMCUwO6N
9f3rHnYBOEICyvvsuzYsP9bM113FSOjpxh0yZ9oybdaCRdMPlM/LvRKd8/o7KzxekfoVYPNeh//W
TgrGFUq9Q/eOozNbsozpYeDPALXJpIMhlmxN390GRMH9foLoYKrSGD1xhTUu8Dr3+41aIFSSv6RM
6C1/kQZP5N1WepMnE2od0XURjZwywhIwkjv/Uq4+2KD6pCbOwXusTkrE8uJfg8FVdWVHNL/8AoeS
Ufv4X/aBK3Qt/T3Ow5J7tSt5p4gEXl2T+qxsjhm8MvRv9Rk3Cc5CvyUI0aRpdCspbR9iEmG1WuNC
wLTNLsmBP9O/UhM314+toTjimcmOhQiZj/+AgsEk+TOOWFEAUZ+2K6pDRoTyi5hEgfobA2seP4Cv
jUWj46LusG23gXhkBo7BVJxsY/c2LcIi86QD9Z55brwIHVO1msmWU7B4j2POj/MZBSMsqK4xKolX
kiG+EPNfL6cSBJACjDyG8UziHHdOPkF0FbRJ4hw2xQcTA94dq2XqDV3Q550jPt6oihnDo23rkS3Z
NPdDAqhMn5DhtL3FT0QzD9/hsyIKW53bcvxYRXC7GVV5CS4zVE1WtLnJZHpB5UG6WMyvR9eybpb3
0BhVHq8pXZjSj1uqA7adWMXWCS9YXSK8lifxVVcdH7Vj2o0/Ocakvj1SLTHgSSAQseyoPPdlOk0h
iUPrCxHnGo65Is1QFeZZQpp+eQdFby47IzrCyU3XmdgsPIjH8knHXeTXpv9I8bQiiqLH8+OVSbq0
YIXZfY/QLqSpGCYyOBxUr0HrTSGCY3ZqBGBfLpRv+HpGORPTMkH52wXVCc7mSeFjarPEQuhbcrV1
xt4s5Zg1dFPP4PTQJkS8gjSSNjDKF9WQRZmTp+CDL5gO4XQAuLFXTtiaHRbftfDmpMH2igzqAvdR
/+RJbt/7liimNPleUQuMo8IDaGRTj4jP+0u0t2AUjgKnVFfSRCcToDd81AX/idjb0yXDeU/QhlM3
iQToGg5jQD2JP8ycENyoytmv/i8LxXGt6oCp+u4vByhKB+MDh5SdcpjU9dz30VY9hbRLan4MBHg2
l+orYNlg85v8lnhM6fkAmplS4k6cPlb+P+m1yzaZPDLsjfFF1WoLYOHX5KYr2MzP+qCw5ZU6lJht
ZaIa6ZKtutbvBN4HcsUUVoIyBUHtWOWLud/SRbvBXkIF+++xeMipXM0YM98NQr15ed3hi96i7UZa
B2HVKDzXLjlW1BEyGXD/b7DwTCVA+A5oxtYFQxh6bT/Jwm2NOzKMmb4/ljaakjR6PpeuSfnjeXsT
9/Jt2/mlSHTXjnDJtSpv39JEqJemz2c4suSo0YcsPxg3JOXKQ9/AYlSL+c+9gW+yE4huuQi9eoXK
0UvVlUi0MgbRM7QvU+glnRAFoYzcKj2HhNRPXSdpMgGnHkSXg4EoCm8RuUdv3CX+4H9GZa4uLACu
wXhh+T2z5Ng5yxEoX3nLr0U0h2BNIT3YeDiqTIcocnpFto62exweaYnzG+vU+TQpIXtE2FMkQlh0
8eghRNgjIn4ArEvkSrr8zBgAQ9G/kPNbEybshkjxFFHsfv0vu4I9ka6vJoM34L7cc5ccqK9SFvRF
Zt3Yb6rnWU9nrZYuarbiFZvp8kVch/l6W4FvRXEPT+MUwxruAAuTYQ0dBvHctwuoircqmP19mr8H
+N5QA2YzBIxJj/2vXKjPmsnPbL9M53FSEPabplPWWKwHhKfVcURMJ7Dn/wxxrT2HrwzSTJBaDyRj
K2Z7JvJwyrXi/TM0Ax3YcvAhTLUTxiFljNTfZNrS4WRLX4RTQGxuFT9mt7qGUAq71eJ/JpNlnkMk
1ZruoJFRy0w2NEf3EehNPwLbw1+2DTBG7DiDIQXXaJgma6g3YH4sS87FG+hX62viZZr04ZhlayD0
iSwvefuK/Ontg7/3+vIHWlSDWs2Ko9kghbeS/HnMJ9yhFcx49C0LA8yhK1LmjWhSc1EJd2fv6xBM
rIeNss95440e20qzNnGX4N4XTnM/6fI8XyCtYIu2jUurA3gxetyAJ2BKvCGBVqnRq9jrjyEpo0rR
Q7mcLYNgVp2DwAM/R9oSFiXWjfKEsaAsrZIOKIbOWwr+RmKjIiubFMMPSZ01AnklZIgw5Far/E1A
RhoiPMdi3hbModQ2ilMFL4iRUOuSeV8I8vL+8YCcZD0THunOprRPPMNoE8LYCMyaRIM3/eLtfzvK
l/LR9y+5iJXjx2nFrATm0QOXkZcaA4fHGBIgqZXeZ6rwHwCW1c3VyZd67KdFgiLOHJKiW1qXA2aL
RkjqgxffAjRv/lMwFAmRlgsA05NZPdJT9RIYGZAwFniHlHZR/mgMeGdvGzsEDJP1NPMG0+/nm3gc
iOfgKbuvuL7m0bb/EANq60K4BXiehy67YH8dc3b7S+41JAJQbXF2FPLawedDZ3W/gd0vI3osru+2
48BwoEBuE4rXfxXNJJGoADzBFIBRTN3fvJR12SwP6AFTENWKI28zYrdSplxNHFXqWv0JdSrgCl3E
i0dCcyO66XaWMA9LeD4E3dWSF/BS5AqGEfrOAZv+4Ap1iup15r1JnoNa6HncrJEthanGiKGRdO9w
vTt+9rikXJJwkx36XjzNZvoFIeqmyDMF7nAN2ENla9JWdO9m+ysY8lnRV1I0hdeDY3A7eOKQHQ1Q
Nx2uQPNr36xhufYK5LJk/Nvw4axHeO2XGKiFGDHKWWWE6ZVp16dVJDFGHbJEIKbP2r/qtxA/snh2
JchAiomaepfN3JUcFXwaRE4GXz/7quC4edsOmEKX5YL2yy1HSXZ9hulplRoC2vmGKE1ydZJRgkc0
HQYUOGTknsKTjfEN9bMzXNkBBH1O7W68XfIpEnnydBuW9wH/cTje4qEKpk1U7b5uf79R/sia7Mja
cKsomkbesL6BDqW7oT+vrnb9mCiWpZOZTg56S/AV4UPQoypw8ck+s3NAG8LXPTfx57TDZiqvC9cJ
Wg6ZPESLfAwxovG2BkZTL+54THBZwBlcRcc31fuQo/uOCVXw38cbzjL5Evu9dIziNYjYDHQLjcew
xZGS4M0m5+1NMR2tnnLMFwEKfSSmO+5WRsrK5vwnfIZ1lN2Dca7935gwRVtJq1ZIOVyhkkp/uxLI
jmo6UjcUfhfdCtkSJO1srqyLqPl+u2aOfnLtBBDYVpcRml1bpcXZZZSSB/2VgCPAV5e+1w4QS/Hx
1j9lbwF3+ihcCAnkSbDcC3AF8LPqq7cnfzLMsQLKN2c3Cj44a/lgi907e0tLoUIXsU+67FNLMxOG
l06O5uAwwTtkU1ghkX0xtWCJMwxwN7pJ2YyEfXXgK2Kk60K6SF8aL7hNdtWs/4bVP1TKIEP5k03W
SJ1jvxj/0rDsCs1sCwTLOb8pphlbu6TAOBjgmD4KNcCda9K9HLS0+aLL+VmFOftfxdQafrEfufqR
dGAb0TcVh8YgLk5ge0QNxFl6ICvkk+n1BiYs/MbO0GojLryvZExyEcLNcrxx43KZGSzWGezDgh36
KOBDFI5TKQESNOo+1/AMiWJRDo7lmxfomWyyAbmEbPr5VCAecjKSH1ib9D3K/m8WFelZfzcJ7ID5
XPkKD19Y2libzbBNxyXo4+E5OTHx56vyrriR0vUF8Br5Aa1ugyO/8UzJruKfy+Aj1sfC1+elzow5
zeky30n3xwRxvwy/4SGahG0BiRfcc4ilcvdvReMkVGttJ2uhyvTjiF+govoyWlsr4vGyLIAwUZM1
NamRoInwyRpqSkKLznINt8ZbQifottDqmamm+eHitjiL8BxUBQX+JmfyXrmGdrLjL3a0+1sNOpcz
Fw7XXDXddIBqArl0k1UcYopvlOvZ3R9b6uIAe/H6wLFYYGy5Yml5TpoToN+jWS74AR27ILZa1RnS
13AEaUgR5Q9vDFgvjE3axSBkLZtB6FNeSR2xNNBZcym0V3I+yDdvZkKLdOlAdmTVvp/Aykosn3d7
bcVqxBY4oCUmfufufhHJSzL2ZpQGT6E/0irub5i4uxtliqRUbkkDe7Gbc/8sGQRg9I9kmq3fJwrM
Mt52/eq2oviLhEOb7RfORqp/5j8x5aiIN/kNIzvDbeD6Jupo7NdRo28yc7PqkVsXaQiA1A/7nEIL
Ecu+uTjes3BLlprv6e+ZHJVInaBx5MLWGgdr2wg88tQfvrQhya1zJqG2ArnM+2XhYy3yrnrcqGtQ
t0OsdJa3Ro5lWNXfEE5B+eaE2RZSzFr1niM/KYRK3qYexC7VM6/l082tu5B7ZX1q3bGS5wctPbt9
lk3zu02lN0kTzLyKz9oeak+yoWtrAVghHBMkEidjulG9scFPa3ibDwwKWvlUJwvLy5nG6Ooqume1
rq0Rzch7VHOrvr+QInTulnESLzAwV4IUoXuHVjT2MJPYC4g5FPNPQ7E+T5baF1q7TMEyQiPyEobW
V26IEIiLB0fQggEfBQXDNVWwa8XOTz4BkLBqCDrrRweYJ+sEEQniU5gCF3ibMdVO00fDK8oBCFaJ
IB7KSZv7Fg4lJKIOfNVPajK/Ri9LkJHldzPTIgLjTusNyB1cwDNnmQ+cvrmmNpYm3Xgr7hYrQP43
nL8CPfemrGJZ1AQijBhCHeGuIm+ibeiLLJefRK0AUzVM0gG9u+Il6YpipM6nIJ+KMrFC9U5Arpi2
DEMNHqV8iW+0c6Dy0zoHxhiv9mUFAEGuqZp1TI9MFunvNJYIHGGmwXB+s5FqkSf3ff+3LQRXLwCA
UqDJGwojWIjpviMNkz5rV7r7pLVsF/TSmLedG1+SaeTKmkw7U695xnVmvqdcZuYYspge0tojlTMj
TDwMLWnCL/jlHNJKR2fmlH6VyKqNbk5rF4qbYgW0OTGqcYFgXSbjl03zNxdZQnCf6mPx05X+qk8w
QYQI1HpTsFBz50h4OxEvris6DPHU+FTzmhct4okRDtdI+k7b/udpxTA8mP3LGQKqcb02Th9044cM
taivsq256R2vwOuo/CApSnY1I8qcv0Y87qoyFG9IfOY9mYDVuToFL7hCpOX25b+5KFJ4wXXoMePu
J9E+8TbGYbOUW5FZhtd520k7SY25eXXWIGFv05bamQAnjblt+t0t5q42q/0u1pwc7APueHS24Q1A
Pj4szZAeC982Pjq+DEXEFcl6vtN+w9TfcXhCZgFF2lxCylCtfw2SOmGwRIguFxtSwCHwkuFP0t0Y
BRschiUCDLgyd6YqA01RPKo9WxLdvMOu6xetYyiq9MFj2QN6po6L11fxR6P4GlO36fqn14HQHg/V
DjhGb7rjpdzMUAv1mss860vbiNJOQSYoUO5L7IuPNfJMoLUDumwS2/g/2swPTjPpOn4oDeZHhRKU
QSr/6MQKSbWsUdIa06hDqXcIEKUHzdNU5v1s+GaQmuMaGzWte8CwWEzw16EnW3KUBNkN2I+QxGkX
CL0FRSCdiZHXdarOU9NhXjaolUY+2f7ZoTehxtghUrmiTrHPRHma/uVQ7j8bjg5m9QN3fwUMgZjv
aAD90Tt8972EMkb90drMFS+BZIbHXP+K67psIR74Xcd6Iism8TlX2RSFlOhhCT6DIYCNVQ0vGEYH
RMi9HMotC2FxCG+kILa2PB/4z2VrkSC8mmFLladlJA6LhEMaaXj4cayLgpigouenSr+laZ4zL8TL
jIx7gMXfzN7srcrUyW6Waf3Zg4JsXQH8smVgiPtEaCKdbVtFrLqLk6/yyCHTzgz62ZzEa61xB/Jh
+A9J8ztKSWRehEbKHiYhblraibS89kecvxXSjCwBSPV81bM8brWwG4uzpU2XTesKKNjSCYrfs3qL
fH6DJAJ9u+BNja9c/4HE5GRBEbpw3aW+VT07qpedE7VWXDV64N9d9zDKBxCyD9IiR0IDT4q38yio
/2Sn/3FBXAAvNDyCH0nch3FCLNiwnp3eEmlZMcDFTw/mKm6nRYQX1BUFbZSR10UX2p+Bf6KR0mCr
VqiUEjNFk1JgK6tjuhwGqXKxMmNpTN12GBAb30F7s0yfdPkRdI3c4MKdoZEigAwBvWFrWcp2NKGr
6bmksWQdqO/VJBX/hdoCc8CSb9KjY6y+au5XOSUCrtboZAZAUP/+wdWFMsG3v1AG9wBY1UlxSWYp
i0WHc9IEpl0RJ1Qn07U9G3vV1BUkHeuiA9mYe2B9zmuEvwo/Ws82T+m+bnT85yJosfUjYXus3vZW
Uv2FVDOiU9i3A9ZeLDyKOVtoXYRqPVb4/eX33bA0Leny0dXwshHxkHFLh7U7p8rIDBCJTsEBt7wg
hA4qhhp6F0p0ogmI+yy9WfwAOgkHaqdA36+7aUOdCkIHuq6SXpU6aa3k1x9Gleg+ar1cFRMtkeGD
2ZpkyqY6MdwYnHsE0f5+Bc7dG0rN1Be8Cry9j+k8h7CDJrXVzUnUNJfsmE8VNouzsFNAMC+Ye/v8
IdLLQGfvI48cLKKBriDM61hzKiDhCjALccbFgkJOd14BmUwevMPTLn2lQTTnjBu/6brVgO1xeW37
TkVA5Iuk2iShMa9JgpRg5ZCx2mmL4eUuUFSE55ThAtt7xU69IXZk8wuuEDP1p1q8HIeIC7XM7mu6
eLUUiAKFNGyuak5wPVZlPTMAcCzte+yP6NnS1ExZdjxE8wpexHg8NvIYL4JOp4C0vRfLV6A+NSHk
6HB46a0/xaHkCtkUe1jdvsM2ePD/v1CySHmmf1pAHs3kT9T767wms2bekJ0J2wWohbATL/RVYx5H
Zahb7R9lveJCyHZfUrE8gZQUSSQXCwDC6ni04GRcm4o2yCxC7DluRh8GfuqJn0CYQ/5vrm0gZ4Fc
SibQEpuVA0XtIhBwtlzGgU1zR430xb1aQXs3oJiT4tlK8wzZB2kzHIWHI2JsgZS3t0e3TLgGCPQi
3YIVFyEgxhchnXw3ihcIP+f14VmD2RbWBqy0XxBKUQfpRNf07RMOUby9FNz01DPTu9uPDYHPRoN+
uE8DWdn68phICbuHd5nMw961yjg535BlrxAu3VaQ/Qo1q0WKuXQesb3jBDU7jceU/d2/DB7IZ50R
xcIBadc+E0gr4LRHVBIPwZOl2ZccyLF/YyD29CgQwyW2tZnYx73Xc27yhh9gV7ANqNSLrI/DmLW3
b6Lgc/iVw8kt7EyqUxv3zEzkcUwSBHmqVozyPlYivW23femZgf3JdIQMDT4UMRrFHti9UaLIvljf
UGUCGIS5aslSxJ9Ro1XUjTupk3PmAmetTUPij4c+Fzh0IJVFvA1+gLAcFWAnuvf2G1hv/Us6xEwq
Tmzdvh9Rapr/TS/mrULluU7NC6YMUue6Q/qrml3d9zeJkLUltDqgCAfVORMgYez/SvZX2p5Dv4Am
kXKlz4hzeFig8OacXYqMMpOtcdQiJz9Mtug7ylU0VHDXxRj6X1OYFpsPtRt1vgbqOoI3ArbxQ5o2
0V65RoRbrnTFma7IjCsGDRCg1rFielfAEA5ERBRWZlDaz0+tepNWmj19Cg4yloFQu0gUta3KYduc
6C5XJtI8IG30vTXxwSX7rNT21lh09CSg5atAjQ5SiA8w1MCxWXQuMNHdzr7w5QhAYRLpk3bc0+UE
Ycq57C3easyNm3NL0H2ronEev7rHn2gQhynvDmFwLEoE8Zd/JymPbutFxWE8oAKC5jV3C0XFpLL6
tY30C6yRqJI0OT1GaaL/QLodWJx5U4nExOTgjj8bHjxltrs2fkZHmvoP54l00LI26wB2VtvvGfRi
f3laxUMleAuoUteCIAzsZT/KNjneGkX3FyoKrIBqHyI5ItGBEggpnWoCOGbK53sAPKq4OTG6BiPq
lfDTHRsByr52WlZifdr29SpOFqD5AsoUZYt6eaJEjWnb+pDe/6/ZJmcF9tQvYSRBKvZMOyGaEgHr
4/5ZOHiEi1P/UXoKdZLduHSUjpGZ1U/UyA1YuPyfI3jNp0F51zim7PoZdvrxH56bpEQnRKU1K8U9
A3vcdbdd5l9FSKQYycluV2PQ7ufHyqVurJz8IpbreiMVfjHHv6mwvd8wNt1piA/cxT0nT5gRQXOK
KSkHturGNkuvZ4aarivev0qrebnKEzNXkJoci+pWjCotneVNv2fl4d4ROVMmH4JnXcxHliCu8B9N
zVmQ880hapKeo30UeSB6xmzM8fv67E5j0ub80hHGMIKiVK3qELbCJ1YvdrhxP/ZIgzJiPIFWrVaq
DxMVAUYtE1+EragQI5kiRGCxBbWw1AUyexCwC/hIfqot74/Gqr66sscOxgt2P0Q0Tzyo+0H7GK4y
7h7Wii2Oh08pop45Nq1AkMNqnXcuCIeFd6ymfhUVHxtcf/bXq5CcrSwR/WEgK6l5ICUfuBOSwNPm
klo1s08I3Koh0fVBLTXsaBersVqcIsHVORqYbF6jBXcwmiZMjVBXk5XfYNyK8Gdt2nfmC0oUhQJn
5wfEqLlMmYmUkatb0PPnVEhQ/JWrirzyBp2a493LuZ/GeYtb+kyPlmLEkF+vn/SNcB7LV5dM1Wo5
3Jln2dlnwLTV6UBNssGkyPLVBp/w+Qto78eN8Im8FlJXusB5u1G3dh3/gISnWApcijfPeDo7YbhK
sjG/rDof9S4WtBk3Ap8chHVziOfyzQNa642HHIGdebj6vmzGd/SHTXHAvYxHRclcbd03oHIfgz+C
x4EQQp9H3ESplMViQtXv8CxZ9WWbslm65ISMtq5eM2IIIAqECrVgt3zrIxPSjwy8YitxHhVL5YTC
S/Q31N5JSKvCJCdln5/ZXmetPSQYUHM0LvseWqUuAUtYms4AQg/3k5umbpUFvzB6WnPSAdn32bOs
DDRzZvzeYHm2/5SxGQu3CPkGJxvDpOe9qw93Kcsd0xvKxR74ld8HyBRqcA3EV9NJCz0Awfd0qaYv
NCs62Yl5t6pc6L/9NGTjU4b+hpaHiB6I0OKw9/CmHe9jvOzGbPjsR8DydIvgndPFFBtS+KNdeO+f
PtbqByAD1BKa5sV0hgoNPLAQfGuiDLMhjnAxgjlDkxWD98+VEXliUApwBBxXgXPkQ6KY54xgXwgM
3Giz0w14FnybzKlVoYqv/o8EPMKTUQ09ZSr6D5iQNp4iBwOJaAmFA7JtZShza6VzHjbLwjN9ZM0m
xs+caqosHaONssfYvDnDSaTt9ZfSI2IK6fPXBYJXr1S1YnlM+B2wBPLT75H3zyvcP8W0jB7U1q2/
eodrTNLWK3zuiUVYeFnYdo/q8Pvg4vR/72oV8uCatjql+6QS8QHQoNjSq9VRMvqq8um585o4pA9b
AukzcWt0SvJa1mbBc4RIZ0DlhU73KJk8W6/rTWxUTgI4AVxRNiJ2JI2XHFJcpcDqu9HwYw8kQZRD
DF0VLCoh38rFCvxKl0DGwdTBmCbKyNpCDR1hGEB9YjAMMEJ0Gh1C8YKTF0g1T2mAgoMDZkvpTN7G
K+tZTyg2EotWQIK79yIMbOEmuffqzzAZamh6O8KdFeQS2obsY3CsU5Lnqxc5hxjmrAmhzAMQmJ0o
9HRMSkpBBt9iuezJrU69HFHDX/N0iZ9jBEqxHzJZke0gkl1+VehOrlPnbLh0GqXdgtGGuU6yYrni
AaEtBe7rzKEkLuDxiCm9S+q06axRtf1ROPhGhwae59Kcljj1ONsX/LBdR0LnwEt7hMfe+I7PQyD9
1EInjWGdXoYqFvTSGxx44Sm0V0YeZmUnwJw3GpxGk4s9ek+A1OyKu5qSjLiW4OAAA7fzdKkxe13f
y0Y8KoLMT4G7bv89Q/9vej5ZNKr8QiutiqwwHxP5U4hSB3/5cJb3qVAmbJ0Wo3RLD6lUeqnhBuFd
mbMD/wXKeKV1EZI+8Y7FXgO24kzDlcvMp9xRzgs+q8uk3UBuCVkxyqcfiu2m/jAQ78YQLIBhmWX1
Q/E4iF23PboHjS1qx3jVw+ZiRxN++DfRgvoDMH4dXne1eqV11IyuLdOBH2o8ccZokHjoh/4p/rSq
dQiz0x+7cGl5xpJLmBQ5jMP7QR9YhidO8pYIh1H9W5IBjHSU7QTkNNNKXbg0cbLAtuLB2tkY2Rjy
KksfrXDdAz6yYwHRZ8kUgdP0elcn4rr/Gmran78T8nRizebeG1fuRYUckxGZk8wbgrknBXTiWpNf
nAxF3pi3qCBtzdP6ZltCb8pBO0w4nwfbkaB1jVkeKW23IZLzo7ZCTuTygz4XYaL/xsoSsRVrg9+e
37iA4ymn664MSGrBdjFpiAtTjSmH6K06mj3lLhOuSTp/FQVGHn8nsAnru1zXD/PMc0T3aziMMJzA
EyZnGDX3r5460tehQFvez90IrPHOPT22jeqA6F+hXzvr/Ylpn6t28w8Qsruj46/W0GIHrVhjhFMk
6skqbq5Wxfyvf5yvpB2haGIFw8ztSg938kX+ptOFbBBBolODp0sUI21oDEfUVZRB025+3t5bD3hU
cnpQ5rLQ+2646CEfCmLmV20nHl8+vhe8UH3R1zICpaJl+k3PbE98Pt+6KqmU94pOg4x34mwHA+mD
h+Vd3MzEyTrTTuh12kvPJP4rWaCP/2lKL+7XrV4Jzslw2kPmyXh3CIhW01x4VNe2mgY2Y9XZbMyj
9A4cpCHiN+2yloSzggBMtFRZOq3bN3I3Lzo59BSDzTViPHg6Y1QwsejQOrlBKoz/mLVNxxdM3Mqd
8CTFAaI+12103txWDO45n4QXiin20hJAV/2zVWfGLdYSVPhXms0YcVCoH5jfu1FmSl7VPDaq4BLB
DX2sfz3G7Wtxl98olTU+RJtC9tsUdxnNUO9zOKqpdvgenraKqQknhTbYyW/OqsDmh/zR6z+8L5BM
6CcEuSxHSM169opN3XOvK4gZ0fTUSZuo4TI1v4YaUr9jjkOY6YGZsR3EK2deOHDgCfX6EqbWj2Al
KjdAkMOjkYq2c3zDfXvsaWIDlq9mg5uiTvwLuqha6kCZ4LOV9TEVrLjEXKtxZIjd+/QqdxcYD5Vq
qYBuwYxMm19QHwjTlOYEh1Cyca/eOG9H6fjpRDgkhXOeFSaRPlYiwCy1TV27e44O34XLohgKGDes
dsTxNff5IO21r28yBvvi389zweVxt9DpFi3mqAb4w79iofzJFOisSBXRZrDm6lG1f60Kga/Ec8r4
N/aekEvYLXK5wOXjGdH09tyDLZH5UANo7vPXg4Z4Ehy5p1iSKGXAJ6c4S+xnGZlEXMFwTFJr5YpK
1DSTahNBRVMqChkZOYDPbG7x8wLLuJ38dpfHXdX3fyoKZIc1mMR8EqMDrGsK0mj2lChkres2l0ny
bPcCZMzJD6K0z14MqGvpVIHerxcRn7KncwZHjyQWYYZPSAPDbAh2Gy5EnZEdvfukgm2DFWtlYEUf
qOkTBLTWZv1SqWvVVuE7YiG4g0np09zTYWL0TI5S6l++MyEUTTwu0+m1Zfpzo6Kns7p0flJ4Ykpg
gnELbUBODhIqb2+d3Sp7dRf1YEfZ+VS/cs2iL8nREK1HbormuhsQddmhwMrZ0xKIZvDbfj9NLE0s
hBRBH5ec79R9e19zWf9vuXhs7G1ePvt0/WqWRI7qGKPdXePYaZsi5xWd4a3899qg00Qt3xI/dOYF
W4HwpgNhPH0FOGDqH2I0rSC/RK2sMFfLsF8rLZW1mQcOWT10XbkyF7/RtE0HWJ6VMfQb9DNSLyrK
jNMjDLEVezQ0PguyPX/g4Rnyf1nMuhd4I31NqhH7V/RineLN2bo3yR/EfMegXx28HgiiFspN8Lr5
+C1B5lVBph6sWeYhdYi/Ztjgz/oTjQ8ebi4ktz8ziiyokLwYzK93v0+6TfLX6cEUE6csAiBxd69J
oK1aGB9QumTQycIawJUGEe34gc+NilT3RZueY88hXL9fl0WgMhNOEuv22H7/KN08+z9bZYM0wwCv
4KZ75rnHCdUAVlohVjFndY7QjAJ3mOV4YEjBP9dZZa1IuFq1PstbGMOAGL4H7jA5n7dS6hJnz62R
XOa9fprHUD7ZJfmXdfJaL78+XkgmM77+nqERLET10p1G23Ey29mw6fMVxqA2jV+HxwAbP7NGdzxW
m51EVTH/JK9/iIShrGfIotadyrfVNWh3l0kWnDDh/hE+hSpJHJJfTpO9d+LUr+/oc0hoaK4/XTnt
zBMMmQQT7VCIu9ePOCo6HeaPnxxMQiFXGK13WuIjz8lR+TvCoy7iEfKxsYNk6uKtcbDr9+Moe8R1
b/B60OYGJgdOTibHH/XpSeeMPFnN0i8X7MOi0NEEYYqe28VB27qBI4+rWzSZ0O0/HGQCHacaIurm
kjgaZRfAo9uiHSn/Vju/3o9wWXc1Fp8fmGwn4WqmKI3UkUc4DvIJnYl39kis9b7lgJPiRP5uF9Dc
Xm+CTx1Sgu/uAcFbpDRqki9sebl3vHhOZxtofIikYBzqxXeunKGhWertKoMDMFdh5OxYU+jDU+u1
2kXcAbSrjPaLcunM9SHUTNBFgfrsi9lVWuDh+EBfdLye6XmEUjVUs+TpXDdR1OBWYaD0V63aa06f
h4QVCepOOUWU4pLD928iCI8p3q1DNcX0QQNnV+fxG9MhCkU5PS8lSfFXazU7hS0LS4cx8YDQM9JK
mmQhDju85d+ykTgK+RcUP4+8+D3U4pBk+UIppGNysaUoUvgkHeXjxJyRgcaynI9FYTZk1a11exUv
yynCWHBScVk1rFuwgcyMSQgFM58PkUIJj6DOYFdfF0zjtHVoGyju5R+5qmx6UzwoCoS26WrXFE8E
wJ3FyhO/6hQ5cdF5IUco0eGKDguRa9KcYMRfJq4beIB8UO1oTdYLD8gpw3kgXp1KptjlB5IYgs/v
FS60G1zBpXr+feE0myAFtDKnkfFQlB/lKcFf+5oGOtZcrZ0Ksycs0wsuJhZKOS/rRcOgUXi83uAt
mLJW/6jQ/Fx5so6DulzzioAVbZu+YjzfUW1wDiSJgOa0XkspURymhcU2DwQ7gRHMRvzSP0VjRRJh
GVXkNlbvLZl4CmFEUtvuwZZpZlBM6IDQLsypRj6CqdNJYYEBeccv90yfp4hazNJkYIgAVvpJr8Rj
1HUpDUDnLUlhXfqj0nou+yIjT+nPnU1K1srCbiPT+SbG6jvdy3KGbZXDtSYCfSS3rbprMKfNezS2
+LXLgVMvs2y0qRef5gEWV1hDqj7Mv59nKVzveFyIwGGIGEeBILbPwVqXdYVEnRzGCy5xe9Z0rZ0/
/yLiqKaEMJsHg601L7DC40JV8qzYGkrGYV05f28lTHGmx60XUQQiw0jyfDag/8KrPTYvJ+nWGcyS
iKJ0KoBOSfAZ+ttCZwPlXxq2YWtgolpzOqqKMoghla3vkXn5Pi/95e+wleIXvT1m7OsYugb4cO5C
JmTpm5GZIO5KLu79gPe5yaojjvj+3YyubuyH+mKtrIok7MLo+DJShe3aSIqu/UG0cA+smYdFsyrA
HKtOlFG5wr1IBX05z1/gL0sYdsyqj3O54R65zmUbHIaWqww0zhOX/N4db7PqN+QeGtyPrh7WqOtC
TkRBf9DEEUEj5UU31U6OjlODbgYLMKVVXossUyAWk0rIwW+R2or6a85m73gVCCd2jU0jU+d4MR/E
OXSDM7MKALvRf6F8bVpKbmTzGknXUrRENaeSAqufO/QivDJngaWudQvWeBR+2zf5P9U2wo9flS04
xbqemUbbIHwRnP7bWcIbnO9FdMTh0C2EcZHnfrghHwVJEcwXMekoGHKjgYNZEJglK56Btg8Q1UqT
N86qAtaiFINu/fD9Vf9ARiABwUll4qt4uFxtCfSvKpMOj9QPL83U2gfWj1l1c1M9zI3dKO9O09Y7
xwc6i5sa33EiYNnUKVCPxFiZA5ZNDJzER7oQWR5pjYUAYUByBaWtzeqjzKwjvihv1VPgvD3NxWbq
tBeTKTyCFtUlYin03DvU/vMef/1RlZPqAZF2GZddOTX1kCBNLzMaJmCNU65R2S0pivMO8DqjtPJ7
Mf6EVFbeKeFMQxn9fNNhdwys4gB/52WglmbBTDavj3Lm6UVTZVz39BBap6Ec36rzi2OCBrN+t6Jf
IJ40E1LRUt52YtRLn8WGo11wi9mvWWYEMnBE7UGibA6KmJ8q5s6zsd0C1AUbzmrbv8H6muaTo9Y4
K0OudqP8EQkeqHB/N5bPZ5zEq0+vJGoQI3k5LY6KziDbZvcbV/QI1xNrZwD+p0+pjAajM8FSehtY
KmC6D9vff2vZTta0ptVyEjZ2+GSNL73QAoz1rIVPv0PPtOh3PVdUHOeKmZLmO8Mu1www0iPeewgM
IVhV892KafelADSViQ2fzzVdEcUWaBp0CzfhNlKbUHjrRtXJfc0+upf/brAzXpQ7xjnqF2FVtT+6
uCNeLsISfH01YkJB+Iz/ASbuw/K9G0gECYIAcoC53lv7BcY1OYVScZLTrgnGBWhkM4/mKxL8qJRZ
czUcWIQIv9vVVm4Tnh7pRW9msIyVyhsfLEDQoGOrgCilY7SFGZ+Cp1NGSTGHaJd/nJEQFzrHuOHb
TexKYms6qOTHl3HHW2DrHDh4Okx6Sdzn23+ej63KNXnza1AFgF3Q1XdTMD62zNC4Rtlv2PQVQGNV
42b8nYGexfIPnrcwDb9P4trZCif+eTCNDtuueO1nGUTy9gs7slzKJXJIIyIoOdGDomAI5MedPOZ6
8/Zp4Hq0t3cHZaMOEbirnVrDqjD+J3JyK1Ma17FpFN5z/hJCqNtTdeGmd35JWnsrrAd2WaX+amiZ
L0rNZ21iURqzo5czE9B7tIOWri3sItH6KFNCxO6C9Wq6FsIo9nXslKDWQTvRxYseJtBSm8Sv7zD3
WITSJo39kNWByJZMvLNPKGOeZddrNwPiFD9cQpo8Lymcr79EqWyh5+m7gycNfzSmNL3IoVfz1aXu
NoCsLyWe6I6RH6vCNNRCBGJLeaKIBm63YSKw7rQsB1BF9Z/mg9LVZP9xzB74Tfla9jQfeRLfvBA2
h9VDJNOhIk2hgLhnyc+P7iKM1xROxMn4R+sz1/6IEfUwuAeZIyhOVjHlQJZcZDnoZR1c+LQVkz6U
Z2lbr7DOWk//c7KkMDNhaclDlOxkooABAgdfsWsyFYJDSZG0ptJi9nEPrwdslBsX/3FxlK6FGau8
HkeUYCEWsuViBw5607ZU5PR6nOT2t77VL4S4yZI/pxTv7GodGvP9o3/gxlfdmuSqjbwrbLLi4yR9
fXTBndVIBkShSHyBooHuYqoEe4z2z4ykT98RBQeRLodlH3IKhF6V0fZDhKEzWk5wp+r5AeZQNCEx
B/PwZZYZf2ydojEglSphx+fbWSgXTWJKVuEOfWwTNrUrUUDuczxkZ1xk39eduF2CcvricbgresQ6
hEMaZkY7rPi6qwY6Ce/LkhOeN21WuXO6+jCPAjvFhqsbrX8b9y/kPN3ydyDKRcITeQiIG1ieDgv7
sENFlG95Ygl75c7P3uqiNzG6otXgA/Pn0xNQvHILe3dd4LHwiCg+kh9jNnXdjB08H0YP+5AwU3pd
+q0UTkVwJvgiy1neut7eHq+tL1KQB9zPc4ets15tYT6owKcYuIvhItMBtzc3Me5COFOD10Tf1qJL
cPQ8LYAnayzg/0emzDPFF6mWcSFoNXuA3q3iZZVRzx6Cbx9To95D7cDsQ6x2Cj+6rxOymaAs+ztu
ZTdbvklVvcgT1BLYxRGBY6dx+O/AL2ta5updBiQmQWT9Nn/ETGjqF/A0xBJQXxnI8skKlQOZZjUH
cqYwo+09wG1JWxRltIxTiHrxk20QkQsaU0mNQkaUivvRVTFlgHBEiTPe/sHntmmod4ItW7UYYpu5
C3gwotHi3xAqQ15mGaGI5VlNUxN0vR5MOpw622c0YkhbwYNPaGm5Dlnh8znV3wn0P4bXZnEnU7Qe
5IHEFMcburkUVn8e6uS1vrWwOM9S+qdPh0e6sDGT2jnHjfIw6FzRcaxXW59jkMliGlw4xv5Ux40/
UMh5KKTuO6HA//6jUkBu8k7SwazMZCbC2Mt3VHh3HMt9Qaqxq+u6CSPL4aJr0tRFJfj0kANmETK7
TY/NAZS3sTe8KEk+TNDnRw5n+2jhQwF1yKOezRBGLfU59TyZ1XrC5QtP0RPTVAFFiHxBrALnC/f+
Il9Et3J+VZZl2eSKQcIARne0qIYZw0kbDHu2dGovECvJpWshothPs3Z6BnkNV+gtQn+tKXetZLUO
3yiOS3vsucSBwJQE3Gvtu+KkSVCYOTYvEL5olUUS/RjiyaX3PZK1ODzfWLOWE+2TdQlI/XhgX7+9
x6fuQJjDszeQORJfsTBWhANnH4i7pXeAdT6z8FjHpPbE4sYamUs9fdGP8AMDJmy2BfihwNF1Q1ru
RntKJfZ3AYaev1Azpv8yK7mMkuox1BY3aNJb6699OGXrqPbOrYFAdXQ4N+te2lslDrcn/RJdi94i
QIvSibWHVI2XaeHHvtR2yRj3JLu4rl1cvW/OeQz8rsnJbnqqoaRLjfXudc4yBuAPQpLYwD13hjX0
33LuTvXHOOFOWS6HEuq1fXnQyTYBe+H53603zk4Q+WTNm2zUA22pjjzhgt3OEmJCdVn5Oq6lswZX
eu3V5I9mXk9aWK+pjxS2W7qYfqUOu5iN8qd2vXyj08Peg7S6lRvy901gppGuqPFxmKg9F+cJHQBJ
QYjdKeu0qxQwvJYhL1v2yfo75uX9TH7hIs48Of5PzzdHewWVK3vd+2JSPDj1UrVjgyaBKJNsR+Kk
YYCCoLc1wfsJng68SNWrwvS7UEBZxZPbwzRjeYdfBkeIVkNuliPeeoUrjhiIctDlp3vVT5lhlIlj
yOHlvY5s+Nx3J6yhleITxnrur0LItYedCCd6LQLKPp3wp9j7VOKJmLPQECNXINXblmgWvFBelQrc
vqyccnpnU6+IVkk6DIW0egQIYkzuBEjja/UeplBi/XyUCLDaB76wgCrSnE/VfMPHmu1MpzMasQhH
whea0Uj4Td+4V9GRXry60AlXrqM+IlalWHonMomrokoFkQGbE1PguZ8d/C+iSo8byV33k/LboCfW
pAKDXl08UCTWAJL0dz3y0w0y+hFQrlBPMNC8awig8fxx3hHd01pip1XJ2cJaA0WslHF7wf7wODYw
4aKOYd4IFbGoNgAoeDHF/Er1emfXvUefxZEDId/gziiGKkflVVJT4tgWhbJ35YaB/zmV7fzVphhr
ui8f8NhYAh14CV3KYCOxsICni0x/Bmh8u9d3FgIEsk+YhmdIJoLO2jxn1+MZWaDqaUACsY2Tt0HI
ubvvE5kJI0b2oqyjPeFvzQWUv6Uv0j9xMTb2/q/AUSkxmdGZTPVF8LLMtoYnctiqY95sv+3LjeSe
qNMq0JKIiL5+qHt+QqexTZN0Hs6g04F5FL4sNMrJQVS4aYjmlPfOoVmMSX0UfQfN3BQDoq0A5k1T
itDQd0MxD7h9PQBADin62iiuG9YTbBVY7qGKUwx1F8WklddbxEY2c7Mu2dyLy/0VIFXvqsZYdEkm
JIk6vPI+kxSxcNF/G9wHClL9DWpGDP533rkJzCCo+i66pb8Tk8dchcU96VSfkujODM4BLT9OZkZG
DfYz+UefXrS5Apwu+Y0T84qaBVAO69TcriARIZ8LubQsTtOPBIhJIpdslZAkB7/i4Fx37/olwuhT
piC/JEn35GcePLZt0ZY1dyelRTsvsjIHlYDwhmUTJissstTvOo16bMOf4gwISdkPBYjhsYgokQOu
foT4Qk+6EObnIyEpQfygNlz/ATiH7SeFLuCTBvlOgrCYCbq88IhbqfTqsY/CxDR+8qvL1O8I6zV/
qaLEj3BDeg9RhUoNbr3nMnGFYh/tYO2TBfWzMhnJox+4k6cubch0atliTVnZPzdxIMtqs9eSCgh0
H67B36PnOz8p5lonDirsbp672t312uG3p7cdq70s6YrZ8TrtrpVB3wBl+d428TSrAarKsA33SPkP
FUCb9pttMBotRm/0PMtR/9P9+nG/NAp0MLIdOHY0LmJZSrqXXyYjoE950E16MVDGC5hcDNaOe8EU
Yv+twBA0uMFGlxWlEnAWcjUbmpWb1AvUSv1+e7GQMAnnMWdhcuMxdS2wzqsAlznCqWgox3x9WTaT
fErko2rYVGd7SfTUcmKH24A8+Wk3pFB+9OsEVa5qehJPEeTtRk8PyH9aM4hOo3vZtJmHp5oieIOO
c70stoHCaycBWA4x+Dcc7thaDPNz0ggbPJkNbpU55TNGFhxK8KFUbModJbe55rZgimnZXj8grgbh
hHfMrHRlYUj/Ros/Jh9+IhXqJ318cZJfm3+1GHZ6HCEPG/nYwlCsEnziPHFVn+z+fbpKM7VbfG2p
VNQuzIXAJ69Ccnifk3JO6CiKNDYGmKJh6seOnNiochsSbcBOYG3eCX1n3IgrTLEp41sO2Cgg2pKA
+jIjY/+9w+tkYMwpp1tT1thdarP4nE7V3cl/LjjHGlcgpWT3VknGRPpNTTPeZ6MuyOFXmTnTAt9o
XGS3P/5JHcy8nTe3NVydg78LeZDGT1fAGdUoPioGvlHJmyh+C74AbHXTisLEt7JOQQ1bSwg/DNEt
6Gxjbq2NpHyPCZFQb2IM+/dT5T3F7Avd6Dsf+EP0gtKMcHCcxixdbx2udKrLQqHzYmgzNVt1r8Gu
ax8Kmok/UFClJzgG39J3COuZTwQaVJBvxIBiGC4tDV8I9b/3n8eD2qtC+KHdQBwVhRaiC7P0dz5U
Wa69whavQAVATKkVfGYbwvpxHBA8xqKeZhJCVCvDQfeuzTwXPx9DViR7IjX614jTJMsUuxPTWaFg
9LXvLaEVb39SsH1YBcVh9P+c/01Hn/bKUgRsEpWSyu0PGVZUZWQThlckE1DHZfPWfH9/AS8IgjTO
r2K0yZSj21yPQlGlzJtzxFiLVMvXaplq/umhGvf5J5ZZIQ7hHo1t2HLBi2eyR75rz7DW4/DWR1bn
1X3ulBj6s1WnZrotiYOF70rZxh4TxtQ=
`protect end_protected
