`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
K68kWqWqPTbVd7RedIrheVnh6mz8vA1/5xsgV1FKnYoJDeCUCMPOHQB3+M31j1AswkwTlwriibmZ
Z0HuSgwJCg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OgpOIJqtRiRVtv4CDJzZ9K4ghSt/uEhN2btTLODteHn9t8TVNglevrMGW/5FJOtSoEWQ2JNY8nxs
g2tUJRAqj8eUoaPK+ARn4f1KpuRcRcIG1Xsl5J5ZoUzeO5nAvHt1JfIoA7fMzMpIMys9HvivdDln
wpn/f3pDwUqbjQa/XhQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hLKoMJfWcQJQZYmVNcM3BGhpPtGrbK6JdxBoAvHLCOiKIuasfRoQ4w1QdIQrQ86Bu/EV5PBrpDmh
IGYEGQewn/0TMN6st3TeeFuQb591yNxMpuhjnr7A2vpdX+hLce9hp7Mn3Uw5RfYp0vv77ZxUfq8P
vsavV4lmbkaMd1xVzlMgrT8WLU9bPS5qVu6X2eQqU8bPOAL3fMrKeCZCzoqw0DDYM3BfmFlZPxup
ni+neDsH1Yd6aDH4oqnbFwukwdE/sfkY8KxuBt1IFQRnVn97OGvrMawvlXakh25IeLGKPNbUp7Iu
KLvgHt74NJwdN7ngIhcNiG6ziVSB5mG42/joeg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l0ngr1ZQywEY8dhvw5BC8L6/aPWrpquU8YoARoclF41ZJFviXGsnSW2jeBHyfYD6EQUW0Bx/a7b1
RjceO68F6QcU38BFy5q51QP8F6h/EygXb477z3aB3vtrh5NfvccB4MVA2NHIi5l25Pja/nyxRk3G
lk/AlGGT4IDLRmuiKNBVG1eWQO65eq8ey3tXl/JazI1acDeg+5POONNhteajalcxrd02LwRlg3VD
FQOnaeOvUTm3wGuyaYcp59flFdIemTlIG6Z3auhYWI4F9DKwTiGjj6ivYkZTIN7uulOiQeqUBmdg
OgaE7tjFIHVY8UgnNjVKGkNEkJ0vhogeUlSS+Q==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
um2kjB2m5WFUWrrJMHi6rTSN36BY3C/DmAu+tIMTXwA0hVU69ZqRJbkR2sro5WdUTSDb9PB5x5sX
r7mvFFNuGj7M6mwgqnX54W1M+ohVUB78sw+f4M3sv6UJ9l9OtU3WgA3pv9qd4vO6FdLK4kh11/yh
uJakZxiDn6gCeCgSKewGafeJvXmnccnMKctMTBdr+LfGgF1rfAaHt0AK5jLjF6RO+nxMUX21lJGR
b7H4Kno/hgAEjRoivGpDpATnQFthzp8Qt273n6XFNNA1bQS6R+/4GEBByzD6jkaKJ6lB4co1VAg4
ycsTWhKm0TUpdg7EVS79wkIkZpATLJ3IEvdQTw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BbrVLSvqXjbmRhJIBXf866PNZFb9Ek5W6Lo0cDXG095ZfRJWeHdhkAIjeWJpEY1rETWvArLM+YEY
haC8iEmTcdZE76N9j+jMmze7UlUq9D2JOGwAlHGF5czqieI3KRNVwm5VXN1pulizGEN/Ff6duC26
RtNGrh1B7UYqwOeLcRU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JN/TVpoSCU+UG08+/UdUOcc5g14BrdXjatEZ+eeFgRwEiplgI4iatEH/zqLlj8NmB18Gy0WlYzUS
Y3cs18Jwh50pWKhAEOMGqbzdIgSmzooiCIOGy+tyxt5o8eBBs8B9uliSQQ2D/YYqpOIeumwS3qUb
de1WTX1iKyTJkrvQJ5UBbLP+szMfVkmqNYgxGFztgy7xFxgwHPiNhvqwAWKf1RK+BpIWn7X5rOV+
iGQ5tj8OhzjlHTo3mmNZgtohemF6eUzgpv9wn6GWM7MFRn7+8dJbzbLCYTH/BKEqvLR0g/Xu0qmL
SELPjDwj7Wra9/LIwej0C8KOZ7MGOeRkaehxFA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14016)
`protect data_block
Hl6HxzyWPgI6QecBFBL9i3jrSk5mG38xjrVSmKJP6HUrrUm3KUpiqAXUQoOcDK9vImK1PrU2pm5C
tQF2A3M1IJsHCINQMGhoIb8GUN5nSHL/WTYU9e1WqpOe6M2ubE42lfVgIAtvFLc5x6JcAAZ4PepF
NNhO7M2w7KzLMdXhP/XX5V+/gXjNUcbVCB8DeOPBaTPixjEvF7GEj7x5IjJcVGnbt0nZ7A5O4x4d
keEAIl2q6mrVl4O8h3FtXkHrSK5KSqB14BfXESUgi7lA8K/yUhE+qYGhV6HmlG7jWDW6QAUHEF63
fck3/N4HC7C0+hLmC8AgD/vaDGqh8fvbmS9xMimUEBqtWtciquzt3SoMstcHxDYyHBAgd4Cpa2Fo
Cz1KYhX1xt9zNXtmf+dbLqvXMmxjunQfn/O6LMq0K+kIx7SCtJfClyRQRX+0dwedi3XSq77cWW2q
xvTD4JIZ17fiTPraWUtyRCCuP+Fts+hSdoIZxhDw+PU5pSRddk5UT7FAvh9k+B9E0s+VDDJApagc
zM9yJ2618/9CtiQNHJvMclMthWHfFhg4PNuFcxXPM3Sx1td/HWCDJavZNPNfomLKk9FWYfUPmzm8
vRHMy3+P9xNYQ303ipyG+v1MO6rUnX1N6llo7DhIB8CjuUau/eJrJg4MQ9mDdeeciGOJ9Y93oZRH
B5IKss3+4ocL1l25V4MTMegbdQusW+5/fD6ftodLuY6TWxmRWHrO+9LeYCPtsbLOJeEfCw7qGFAV
pjTLsBxoaxvvkgoVVQZxJhQUGv1Gd2hhcsKgyor4G2zrnH+6NK+glsbM7jA+Q9W/sfNcguYL2s3n
Y4isNYk6HlVzkoGbuUKBNCvSwyr+KxZpOwM/s+9L+exQxwrZ1RzwZhAP95ozEYd+KTIIkgdASjaA
1QNzeJJuK6OeU38GRPtX4jPe1YIuBXCtJodWAFwPTztz/9BHkuaZ1C8pJQNucW6aS/7zVDzAT2tf
sPqgoSzmHMErQQGNr3oNxfL4s6Zr+SOAD5zTH8HXv4QAPgYK+0TN8nQV3odQul2LKyQevSsFsLk5
o5bJbFPKjZd7HXNQNBACryx2SE5eD3k67hwtvoKlPfvjvZ3NfarR7dvoAumX5kF/eD3Q4PgQBs9D
5wLsOUMolYwUpBOD6dzkzqMKv+gv0eZS/2Qme/F+BsJm/ny+6RCGeVHtU/PZnyxT7UD0/CY4Sxw+
VFKzc+Ic7QjOWVph/KlvCejFhDjCYj42kiN/7BafzvMAFofwytCBwBDgAi1D2oAW8O/+ObMER7Hp
beujR4HFhiSG5UNbOZ0qjj+nEf9OtFGNC7i2+zNQXjiQyCy7a15Z0OgLVqR5h1g+qX8zm+9WIU4J
7FcuwkQ27YDvj+LpCWNsAo7HV0SvoHYdjNts5M89vFX69+Ctc82qkNcq3LH22Yttj9KOBjhRnJkG
ALuLQ9JpeaGlbdK0tyGEbNw3/w1X98IwXZ1qxRZfb/FFzk2w7svb8BEE7nkV+zc5rjxhM8uZgrob
z3JfPpOF9eJK+8r09niBdzmeClw3I9bBLaebojBVd7/0Z0pj5/2WRst7c7N9jZOU2xT/f5gcktiN
uNkMisxBwLBUmKlC/t9TdpPadob5ZGEmg8QfKycVk3QVnzAWAX8FfcX1Xjt+XexboZduMsnaF6Oa
7BrP7aUmHETYJIJM35Ql8g7VgcSuxwyf6wuhiTf4fbC8UO8rVgThW4UJSD5G/uMrx30FUP5lKQxV
fJbAzGIogiHWI67S/T9etqxW79KQ4OO3SLirtdm/x/VZUaJKviFfEY+B2cP4ZYaNZO23nS60knK8
sMjk+PeXQv6Zt42Fem/ughdl7XQxwU7rExaQt5j7vTbbTy69QlpcnytjXGbe9M2Jk1WIvKK5oKvd
jxlC3yIU68NDwXl6z8E4prgf5L6fbX0yK5DGHnvlBG2CVZpH4ql40+vbr+GX2IA4iMjMF4ChvRyC
oQRcGzTaeuwpTe7Us/uvVi4r2zXx9PPLJRwrygeEqcq1Yz8YPKZ6CDLDSdQZwSFCmC2cTMIbQ6JU
hgzY3mzVcSc1iVKNWgVIPgk1cSsBOhlYXRBmT1KDgQerMhAdEFkmcVhmxU768xtyGoLssj+w3R6+
O/HNIWcwPyWhHEwsIMpyQaxhPWxdQXMqiD+44L0xShCfjoIoJhZnf2ca47rFjKbkyNPE5orm5jMe
LApSh9jj1VBKSerO23ASkwXxQXnhsUC82XEDAWbXQtqKWRNrhqq/ueYqp+z7l3izxf6pbC0VWhnD
PHWrfJQcBjFry+lKwqR4718J8HhK6sllIF1ORvOvDUV9UcPOnDXwBxJxhjhoapC1JUmFTH+53+sg
oWOR6dcK6Yxc/3KmdfKcX7+plto06Yl4U+SrZWtifg8htyvJi6epMjd5HrriCwpmMUqiOOkxvsUY
iXEoQ86j0y+G6sYHhhR9uHacQzxsQy0b1XsVN/5w6b4vpunKLpkuwNLczgBaMk591Tg/ck5NwMdg
8gsh4Q3TIsu67hDx3DoTpZJMBv0Y2qrqkE3Rx76HnXOLcVRhg3Aklv9Nvu0QWTCEsyEnFnodlnRn
QgRT0VOaAYskKDX6FQ0B7W5uOl2IgMId8CUY80F6kCug0wP+oOYwCbAz5oYiRtJ7t/upeoL3qb35
wYJJGn6VHIskeMqDrpPZNpQ1xW1S02qiIqBSPp4giveZN2eeGEuBQFIAL2puL4V8hf3syyi4zJHD
x1z6Z6aQTFXE252sCdjw1xH7GiE+3mot1HRIm5EdEk8S6zwpK+jjnSB2PLNmfPgGKOtVyxnWPtd6
eyJpLymu+LR+UXSODp6yjljgfuhMRTd9IpGZSiOJzJA/Fy63/TRWuniBkd4sC2/OdEfGdqSsjb7J
NmOxsRhi+gbT0k9ohCBzPIYUpcgr//vQy98RyzzgiB1R6/WquoH7A7vWBQXL3Q/jSOrNdrDwXaww
o3WCTzrXJV3S/UL5yHi6EKoPrOC/tQsVyW++qSmst/R21jc8HlRIGNUQFW6E3xRl53fN7hd1sOxO
YCzt23jJOuZ/Qs/CcCqJZVQD01I3LcpGQpEy1qU4BsoJCHJKCTd/CrOaqce7xXNK4yccMCLNEj30
RFCuil6cYDvtPe+jfXE0QTCTk7MVR7SqI2TJGRgsA4N/+VXtTKxyhJ5Q1uU2cIBfTde5ktTKqpN+
MbOOXPED4ucQlBAI+rYLaZ8aKLPp3N8J9/OoqGuY01dSGPmaPSKu+NqVhvpTUFBwgnzhLupByV1t
wUjfhTrLxh3OzFSiwYo0CSgxqnDmL9vGekbpU+6MG03lKWb9fAY8kQMkNzbCEzrJOA5E+UmJKPV1
ZxPBKcA1l5o8je1/qWFHEcs+jB3HtHYFSP4nFzJ6kBvfGL15IQP7pVSHrkRIsssAeXNQE9InZngp
TKdqJSi1tpkbV7OC5Ny5dQyn9gZqSqUo8lQMl1w7l3a2nRQV7uAbeQjapRGKPsZ1qag0fLUBcOAm
pyKTcMhwh3uS80CNYG+tdsH64r5UV4buT5Xn5Ha6ehX0+VeAxn2PqgJN47mAcubZigdRbdYpubFO
FZSoslT8Ib1U31bfR/jDZ3YfUJegZXuKclY6cQjhV9RclPSVXlLfJ7B1d4izmqvTwDz/f0MlWrQU
1/5o3oOEkXd29q8izfLRF2Ybnaej0eraHxi1DcXkIxNDi/yu88qcHLZ8dLpCzxXwq/3ZmOpmJCPx
768QeYR7wwFDyYGh9ZpgE3WUboMf65SwFxhKnjT12omtuG7uGqT+J8A3dQvVF0kCK2clCUzPeIY7
dNJt8Ow2bTrikxyMj8ymHkhkHgh4a9l+XIHaouj3yfi0Pqj6Jg2y23n8/aoB1PX5AtqU5MRSwrlE
Wa94JswPVvNvfL10T3/XPH7Pp9qoykjIuSq0ozL2i2Wqqm/eFAXycA+PA/QPT8ffpCHAgDN93/Vb
IXV9cO3yvXQaNyPqrhhQDN9mGES5cW28q5bSEUFZUjOzr9bspySxty0UVLi1o8cR9x3jOve8coix
gO5GiTKwOKbQMxbYtsodvwJbPlWJd8/im2/STxv2MaHVDq9aKmgLU8t7Vj+Hz+p1ipIg2lXHzl3o
8+diZOXnP3Am9PnxvdmPH1pc5B9jOMoGwbHgQ1FoZglw0EpGItBwneTZ0DA83CPE/zdJ10p0rPt/
5SXHfRfy076vJNLveVFT3B9J/qJkPj8NJGRuZ8nHCL4C2QX8L9EsLZs/rCyGlT0ZGQHfN4U6i+Xk
66+D5jNAueu0hQaTv+071w3PIL4lMybegwm+9C5Oapxeblh0fvgK6V+TymRThVrxtOiCuxTyOVu3
ZJgQ9kA6L+mCHQms1JmB8+HiOloOdRfvqBGODK+DV74Cq1iVHJtyQ5HP9SHtoghE8JGroES4mzc1
Flc1fZtuLZUEAKCjYp1jRgNqChi4llVYCBCr22enyt6s94K+lNutvXYdDqja+9kFmalPDRK9PVBD
rh3S8JouhlhNXVjUavc+pavOVtjED91T/LblQHGArl84tU8HvDZzeSEODTzcUEivXjJnGLT3xpfY
Kmx1zkScySxfHweCgGfa9PI5YCHe6d+gekEYrh1up6Hec7YdQ9/uUfoP+ce7J3xkVFajDfz/L39e
p9PPdRj0A90C12tYi2MqsWuVfIWTZjKFwh6Ck1oJhrYLlnihqHmCt6Ux6He/Dw8PK+qrRcD/Zm/+
+KD9xHVPh7ebm0iH1Z/gk3nbtPO7R1HyQBBagF7xUfE6bYQ/4BUXaLBSEs/Yw5fInikdyrCGqrSc
/1k4ZcqvInBPYK0hUyRvJU6G6PrgFzzx+0DO7ie+tnUJlDD+aoQrEJbkgK7MRdyaHhaPJf4hRgwq
LSHcy14q6rsFkaOdfeHdB6RWkOaXMY+van2YR/1SAxFCq+KdBWPNEGk/4/MlgeeEQG251ztdFiw5
lTcl+ppwdAjM8xKSbX377rs7YOEaIIrpxNWFTzEutMNr0TUYoEYyA3OtUAVQ8evEfc0kDmgaze/M
hLKJSI35GxYZKtyZ27SFyhLeMUKcgVnGUkLupsQKKXjnCaxbzmOYZP6rYDrPpzZBuZwzF5fdtd09
qeT3m6h+fXSfqWvieX8yM4NQ78iKRvOtAZwCAu2mgercTuxaAQ+TIz3pLCIOO58IVLsoFj6Hmd2J
tFWhXlINqGvdv5CSRT472gXgP/W467x+x8GoGOhdS+RO7Uovo/KcJF4XzQoInEmEW8yDh6qhwFLB
ejopjEIp9selygb7Zq1iCD7pljEbdG6RH2oQHAtJeoU34G/fXNu43n/5JMYq8EFalvLdYvT3wjc/
cQRq1yxdZ2YI10yp28/u3KndjhmljCgkk8w/LmHqqesCglCj3DViJiynwGchWEo4vGLLYDtLTAhL
DCEBciI8QeGivtgmyLw1R8loCjKWsfiuXHzOhEKps7rdehYUorhN3Btqp4nxwRhjtgHqSHQnKefM
z6GjqP3EJuG7Y2snmHtMnocG8P1qrpAa6XpwS6QcjJfi4nzxlmGWL3qqYGDLFGLa7bWFHXgNI66o
5QGrACNA2IeqH/yH2HiVHnv8BF8Lo/EuKXh/J68Tg26T4r+ZJ1dQflOSr35n/Tgh8VT6W5Eli4fW
TMDF8iLdfyiZxAuYTfbRxF2ZBy4nA64OkOWKaDIDt4D/z8wA4gsNDlAqapuJFuZ/6OF/oiCOCLbp
2Hi3FPUc2VGqwMoSt94ls9L3JyQkIBwcXb5humTsaX1V2iWBE1WQsykd4nQMCCKuht/Bb1VccOdX
avzkTpya2fzKb8RBNqwP62XuBg1/+0bp6EtblZ7E9mdr9iQKyG9QxxmZ5ndUlP9W3pUSX3VrvLue
WaAJD0HSa/qRYYXf4/N5Pd2DcbuqRpQlVUVk7FVQhNDjdZHd4XMrQnlyTwS/D/9BPG0cLuwCsVrd
AzkrVq+OpC+V3Mpk8hhxgfHDFR6RE7FnYWvbOjUKZsM8rbauGb/FRZcgEHbCgNVSHpCdfLetXa9s
u2ruW6fHg4d7DyzyGuNGNMh08xVIjxr/aIi94JfIyMZIkaV56j02buRXks23a+fh0rYUBSBGi1b0
R6lYCnsGEuajuYMeOZjF3s462Kh8EXvbPJSXbCbVMS8Jo823MY390PFatd+HdzSI65XxRjfZXn1o
hlhAgURbBfbSRAfa2lFWtD90MLMURBKX2U+RGDd9mqGF/2qZzMUak1pJChB3o8K9YCU8Vj984cEs
/eIB7oQ3R1kHJLMrmZTORsRvlP/2YIZ1OhACjXxTqSvtAV8V6KI6nJZndOVQubNHFp6on/QXI494
+klHR9yFZUkX3/G1spNgLr0y3jW5Ze0oi4D9IXr8cDfzjhNFCcbVQdEsfYyKDbWh6mZ8GbK0vvFe
bezE/q44alwy0aHXk6Hbecr6CO1BWuSlpoAhL5JBsMzG5/Ah/aJ2r7t8jGPyAwqvBqDEb9uGuczY
mVhJyhOy7rfuzDFQ+cMzPCBVuanRHiPrQVVSft4n/PTutiLPd/eBZrsWU6DcYVzEy+e2aWPfdp67
FEgyCigaGzNQXMDfkIHa8wTSQrMqU1bnoa2Ckq9fHMyeBYT6TTUCXW49tYopjOzpMgvfM+9H8s3N
iKn9MgoBGRKrOdIEiU5DZvzVWQ6h8NXFrQt3uljuD4oD+tLPapwK/stmckZHMDoxW9eiifzrJNoO
zT/Gki7p30wxnfvAIGAAOXQfgkyEIwIQYqoIdXfTdQCLFG2R5HiVoGoybKREQgzPyY+G4sDTUoyw
hykSv5psYtzvVTa+BPPfpFlz7c+150+dJR4qnf9W7hBo83IrF4IFnvUiWLcSX7MjK5X5MmXsMj0y
maVPQECPKHAn+QE+6M5Oc+/WDnZn1s2d3wp3pozXzFBl1SB748Bz4zLwxgY9P8LlBjM+j9hW6D+x
5JSZHHAExuv8pJRShhjs62Egc0polqIlzeTA0UFVzyQkin/ZOQ18fFM32iEZkKJcocEENhjSsm3Z
c1i195CGVFjHKoJbK+sRMoDFnPsD4fO4RzLyJZV5e3neppMa0VuboVRtJylYvKjpm2/vs9KwAmT+
iCD0v4Z2Gq21sM719vx/3Brv9koZDCBh1YTGDB9ZvhPmsJ9wMaE3SZtdTvwaOG8d88WPPvxZA26D
MsaqSLkYkcTKQTDG5oYL+VqZEcPQAltZdFw97sAwNChiJ+EicOA0XPklm5V9niWkwjBtLocul77F
fxhEmjircHRejmrQCo24qfgB8O6LN8H4HkvAG6h8/6gzaRA4jJOZ7bgds3fj6GUZD1ChVyWs8+Yp
/dABlO3IoViCuGu6KBJ/9Yu3uUejgQDodJ/gHs+tdNFJl/vG7ghRuoFHTD29cl4/u7YeZRENLtLi
7VAa2I5HF5lhDPwaltV17Af09jFwSYJHoNo7tUWu/NnbvAMVJavghnbqzE03j4VXSmzJL1FL8tKo
RKFk71fYfKVOSb9ih2vGSpF4CfReMBswMDx/TF0Si4HD35R05i7Rvh/K1/4WSFDgivnXMkmVe5Yl
gSeDZTx4Od9qzJrm1rthEH5s4qjhtg+780og7dwgEfrMB2gDt5iZysBuvDzOfMmzJz+Lm6N6yOej
mfkhy+jKu6pOz+Eh5xscxp8jDEX/1RrKRyvqC3KyC5R9PqVGmk/2G6tmai8rJlgNPd5MnB15UBaT
St+DCb2LIatRmqfz0vaAcD+adgvnPnFupHLSnXeK2ZbLgc7fhDuQ6q7n00nDo2H9bR8aHKLEzzvX
CNGJdovljSeYabUdlmJYgScf3pom0/fs2yP0lfv34QpCtaq5su3enHgnWePKovI6qVd8/GzIvGi9
QG2mA2UTYPIoQJPCB/9HzFnFse0BSj1VCL7WNyfW8d4YznwYPG8oFLUFYL5VjceTYDnAyYunOcYe
jtnJO3oOgwCvV6mhwHi2hDLc/8fP+u/6QfCKO/kiMzHiHNTay55m/bLlBoy04MPB229WiTEDaqWR
0LikzpmZiK3EgCR8riBz9i9J8UR30ukafEs3dvCScvaimi/SFlNgj62lJAc8LJpROaB6Aib+OoO3
9FSCq/FOoA1PPXVjCJ+17W20+y/uvB6tNTJ5Gk95y94ZCmdyBXOKk3qG80O2ai17Z3qdNlIVGQW/
tzc+LepAxJfeuofIkx/XjWuaVyjTEQFeguSsbsDI8vS9ikpgOMoJQ5YbA3iA3+wP/97KIUGKyjP2
NT+W9aVxRpUtOvASWb3LMIRBsJfAS71Fw2nBWqWaW5UNoJaHp5+3QPX73cjerjE3sc6SIo9IuvGy
FgKwau75QRlUdSiwPUKO7HOVbm8BARoBe2wCIbk94LoCLKrkt+ooEBvV2Gb6UuO220V16Y8paJBT
iJjo6dCPu6uHlJI+h1TUKCg4rBVnKjSB/qRdM+DRw8y6PltFYrQhEl+argadGnHi1wJDGedzCola
qgakAQcQ1S1BJ0VtB89eRZ0Gs13QUGrhvSwwQwbktw82COts4DxWgbvqN8tWoSgnvBzZ74bLSSDG
LtW1L2pFYolgCh3TbCKOyeJixMeQrZ0/5S9IlcoIapWoH2jOa+0oEUs0szCcrvlWafqITlICjxdL
7CKNFDr1uF4c+Anou0s4fHVSi7E7NiK70KXCOB1N8JHxQoQwrsDTrtBu9DhGSKs9OaFsBRJjPFkH
mDYcmX2DzMjAdfnUn1X04dhNpwLlv92fIH1RPWwXE15tsH79EnDlF+iw8Gzboa4p/HRyTzrtzm0u
GiApVN8wI8dM8+/FtZuuE/3ntTurffm9UAsYEcUkT80DJy145Cj/JqKBytXW+sDOe03XMQbOi9AO
V+BHZpHHq8so1DVUVEkvgLfoc95p7TKmFYZ401f66etB066u+wvnt8d4zL/IeD7PGeBGscfq0yAT
ybJju9LBDdpNmSGDj9n1LcRk2Z3TdzLa7QZCZYh0JRELq7vA8EaJLxYYitQptKAzW+qGar/TDUpa
6UizwLmPa3aldieSamCZR9CTfrXgfwJcLlHnA073+cGYKtNWI4tP1KWSqKqqwnjIQKh6ftsf8FDi
G+FeBnXXj4XJb0AnmLTPTowJirEukaGgBKYJylNyPbTb4LC1udUAq8xpqtWu889uNZhFpFIew3aJ
ut26c0qyceG/l70a0MaMoRXWkrEdpBb87BiS5V7Flb39B7nQwbS1RQOJWucknC7D5mpsKGkFC8TV
aYMnuFWu3VVeJuf3WxDHgFBgHMeQKIdvHRJQctlaSgWgKsIUEF2RimszLoFG2CTnJbbC1joNNKTK
RCLNlcBRtph3fPrIOvaLmCPlWlY6iodg93S46Hll1fkCU9qgaA/5Rp4KF/zfqoDcOLcb1cpRci5m
0nt3E6gJsArzZ46Sk5uJWlOUNBGuLlTsYuN3GYELI27pquWHu6VEJh7Y/kUmU14xpn8v/jtI6e9w
Oxf8cZxHeOVo6JxNnqnWfv+e24y/wnjkrQRLiFv5vNliGlKVuY6wpnWarloO6Ves2uPkae9x55yr
3BqBDljzujzQs5Y+xkEDIz843TV6FybOnSpAewTDnsuE9/i4maDiVQsZVhiMgDQBOLI5nOpcQxZS
DzeRzmKlCe9rYCuWXAUP9QKeolO4bbCsK1To4JnFAw2cv2onCXquUD5XPMkl50hkYlecFCD/JBcD
9DfRlE5UWUx0kIwKp9ZtSSOjynD36x/OAb4WQgNKfFgqjsMDjV+Yo9qIDMP8GnmbdrC5yHUfzDoU
uytNwXQInepvoEAeLJGTEZT6OSGcMOafAxstsrj9Z+/ECVWO0eBF7kZHn6gDK9lnvwRHpC/7oaTY
aaq/PFZZFh5+oOE+9whM+EAAXMrAp6klnBlMSTDYifwQzw574glp1laSlou9yyEB2o5vgMpJDDHM
gy7Tpjtl8H4vnw1RHox+xhv9Lyr0PswtE4Tgw7H7rxBMxU50cNylP14Y0JHY9pkHzOvYPqdAVGAG
GrHDUNFGsqu5y6DSoTlkOA6tLGvj8oHXRq+7p00XodYZN8BkKOlqIyPgMPi7fzIoN2NQXqm+V9Ir
xcPal9OhTcwBL/hN9MuzUM4i06Y8m93tnWDYMSTGl21gKEVzKPFoc3g2sFGzubobz/pb3W09bK+v
ANpEFTkFuTlqyJFy/TYGxRbJ1cP83WKLAf8/11AwnzzPWwP4Z5l9ZE++lowuWztffqa2BxUVDZ6r
tpFbgGtDRnQJpnUeE4vbARsc+UvtxHktaudv3CVO8il9RAzuhAEM/H0w6xRBRBJgBPCyTQ3wN/aQ
gDZ2i/I2yXWTZH2OvDKL1THBdaXLfSwCz8ioqB6gzJ1d4iuemdybDadp7YUKKjVhdBKOKke9S6+x
ImW/lDJD2shwZdviykYPGO3C2iLYHUR3uv6bA8f1zsJQa+fPeX9V/j/3IHT1rXbtxJiY3k62k9Qu
He4IMUfWkzxuWo/+cMokwRhUvDf4iaVZgWCxnZi7WBGF9S57jspxSh7ZNdi3hmDtwHGRuJ9jKMMI
avDRsmv3E1JYS8JqmzC15BMy9Ufe38HL6PLSE9akAaywHUgTizS3C92FBSu8ZuiGQNLPW5xnpCdo
fuzsLIuwowWGvSRywKcSaVEzJoNCD77nwlvx+yFHFhpcaKUd79m5VjL/IY8znh1FeIl7Q/iaMn9i
9wiyqPDtcZDdIWrJj0LeP402Nx1KfN1qK/Gn3+8DJHsfxVS8g3Lpldvg2bJ7xlKdaT8nAaL0ygAv
WdRgZboEbvUdpqSEpz3FZQQ0c0gJjY6pFwZnbzPFIS3x0yqtFheLGvPhzQh+xGntBaZ+EWN/FeuP
UKw8SYwI/eHaclWWHyYQI90nkFGaMZQ6H+4WlA0lNXN6X8nD+iL4cZODcmybtqZsLUb5WEu+nazx
/75Ih5QB8m/rXrLGq9mu4LUSlAJeGX3nJZsjuRmW66YVegqWoqx2GuvH2ov84Vm69Kd87FOfS5qM
m2fhUeNkDMH/TLsqKTA1zd7UITIzW9QtaN8ZvrkzsBEP2taytVythVoZcLE0X6OhbN5vdCKjzRYG
IFVgRXOMYcQ3DF6/VWwt3cTJgI6byM3kpoZRALpL8Nl2vIRgdoF4CzMJKbFC9Wc/PEHDXvg+0yJT
WrdEU5+VbMt0dTuvf3YdCx8uNeZq/o7Bt3kFz5YfVaNXvEH6rb9sKGeKzW2E2mfN2D+mlFRaGLFj
RUXgvPzBGYgtn6hMXhXPLEUjLkMqB/4FF/x0IRMZcGpIrTVqZ9kKUkXBNB8s1eCmbvrGnJt3NBhP
CxCwmAg4led8AyhBw+UjTYhScTBmCw3klWm4f9fNsNdyR70y3Ji1yHXtrv5QyUlR54LU/BylsKPp
5+RruFn2I3OPBA/H2+80uNH0zI3T0YgiYxRqYGbSZW9bmj8xRuWf9T+D3bXMaoV/8LwIGfbLlrRo
bqktNhlfbi/sNkcypZh+YycLmYsnS59NtAPQ9uHLoiSTezEMbymkQJv51Ar5hXECiuJ/+Sh8HCqZ
EBuNGPcyKcQo6cjlSCFIOKcLUM+CL8dvqTOxJuAAta1edFgQxduCBzUqVNaTvmX9JN7E/f/cL7mA
0sSfRofk/qHWSKdOBU/HL8mE2FrIMNELos11ErIJh/T9MaixFdakaxtc9nEHVYNuTS4HmMrhshWI
GPz9LLuCiq8PgqTmCsSe+H+7SeWA5mDDX+A9n9m6QWusYoElGwaRU6H0erOVcjdsNb0IiGGCy/1i
gbZuIL+zFwq+/CLbC1n4zYnb37Xz+o0HrQPVRKKS/BSpMsNVkpLNedNoLZeZKJEKrNw0jEbftrhp
4qbQqT8zAriEag5zdtHrXCFoEnFV2iMK5nDsa06PLuSv1EI2jRLofyEhA/7ayJQV+sp7CoWGcWCc
bbPcAANKfCUPSvZ+GywXB5kcOeiHs2yJlvRuH1kbVpCj/PeTcEf9v8vU88smGgFa4UlMVarle8Fs
vNgKmes1k+QVW1uygZnwm7e2eAx/BD9ZXG+89Sgj+lDzYVinMM8ScQzqUtcB8lOIeu+zVA0GdRFQ
za2uf5RwJsR2V/Q+RUb8wpR41eA9LvsNpagUnKx/E8HkJnMLHPZe0EyevLFKYihGp8olcGRqSZMX
HEqNx1xjIgsKQc8GVhs5HcKVKU4e+UgifRf8066CQZRfPHEsnvXXTVpTUaMOChoW+PD4Z7VJnGPf
qu293z4/rfFZU3U3QW7ztFpnZln5Vjc9FaDoVccwUCoZR9vNh75q4vc8ReoT0AG2smJZycjwt9Td
F85W0Xytmrm+z7SbYKazQj5k1XhSo10UBQxxcmjJs+S2RyI8ZwGrMZsVxDwevMaSY133DIW26il4
12TVTvPx4u3bqiSOh/Tx+isN2PWgzMRAckOnFM8d/gFxp2N192WMvC8bxb1sNC2LewsizxfV3O+D
w2noeR0LEeTLU4mZEaR2qsL9zUiwB5c+WvCHEIpOECO3jT8Namwv+9henkv4LB4OqqA+8bMLnVJt
hGwfFJohRdciLq64is2ff1aMhRJLRxHic5MTGCl5y9iTS4PGD9eVDi+J9Qi45GmOUX8eFdDqP4QB
fnQUXcmublk8i6uDxjKf8Tsfz0vmBBb6Us6fnVtN+cGS6sIPpxPKN+RFztE5ygmY31CyuYheCctd
rzhbfpA4Uqds+yRADJP0OoHHOFa7Wi9g0dIrK5hve0Lqdkqx7lPECTUAK0HmcKSxei7AOYQVCyHP
tHT52XE9rV7A8vlL2m0PF9BfkPydkso8nGsvstQupEAJthmdvv+YEOuxMLzdoN7sf5rJYYLDKuVt
7aRCvqJKxeML4EWkCQtkI/0ZTuVHVpP40MAkUXVxNdnkhcb0OP1TBtiwOtQWIhzyMWV/RpwG5c7Z
/psYuthsB0RIFOXyNvoa/kVzrW3K+MeC5ECFa/H+wpukHq1UmNTG9ZQy/XjsLEq/+es/tw+9+73h
5GoQ2gvjPowDbnnnLL+3kvcjgM+79VSWrc6gh4cC1z66vsuIudXG3fNU2HhvDhOmJBcjWAVpUJkX
ArpSdINP0EtViQrlKecnoDwYs14AsIouBTsTUb2QhuH2hOPmoYb53afnKgirhjf3X1RTDMFd5Qd/
l171G3REYO3CDWFNNXUKb+zg08AD1NfJt6Uj1m3bs+y5Bs0085T0Nicr88CZqLROtQw3WsfVMXpA
3U3d5n+Stg3WO4pmPXKlAT8IdBO0iST8e31ArWIx8T0IbV2vqYailyCtvTq0rXx353ZUorCrTD1K
xONXDfSoTCVpPC3fNj5hDfnA5ALCCwlZJ+DgXiXcs06p77J1wQBl+8JHrGLX9alpbwbEfuBPp0N5
wqZf0YzWr1YpFRk4v7XFUbtQHtjVdn56i01YVP8/IDI8JRF8tjo3oAPAsAh/WUI1et8scvIz1LJp
cWUuZkKZhqKRI2UWvGkX8WCpVBxtzmW+PKkmqa/PcfuvgWAo3FZAtcdkWYfBs4mjkeau6po5k6MU
/tc7RLWHU431ViK6jyWj3G8B4LR/+X+zv8VnxvF5kYyKKbWhOkrAcVM+LmJ1qrf+feOziWKEvjYS
h5p+sNJlZghCZSqb2PGKuGFpF/zejobR0vxzXXBaY3pX2cd8el/4zFX2eQRQFsZtSHyaFixpdnMI
/w2/L8cIo8ycnwQspu8cng99FYu+2oi5VQgVOVFzD/mcyOog/Zlxbu9ez+WCvHDIvi5SFzJrAyGi
GFg4s8KmWXNnVUUq4sdJjym3KvcaOPOeEuCfwcmGQp051NaIjARROlohkcem5M8wCjQM9SnrFGox
MWf2U+YG8bYrzxWwndOAjv3O+sTW1U+xKYqN6KX162/MElbUntlUFPNPqKQpnAb2jg0RVUfNjm3q
o5ZftXeVp7/KtrISd/RRFeMoFe5s3SZuNfJFiTl2suQOHfyAZQPBk43tSCYvvuyv7VOODA5TBwpg
uKGoDb5l02AJve/gs8EksR5D+r8lyuRAFWWoxQJOMDD6vU50pzWfk44bkFL9ygvtbZcYrm4DIuVT
qpFX5d6DY5Mv4ivF2cwzAgAGM9b/fukL7M0nV1BQInOO5701nXka42wH9+h5wfZqu1SrRY67KA36
+qAYa/+nDLkQgkbRowYiFcEFmKXswXQdU38p12uDKJNCoishjZRAGlHVdyjw+2buwkJV6QqHLnnh
/fB4mPFH/9bQJVQrq+KUwxRwtCa5/lghj+8J6kiYiyC53msiVHUMgg7gZ8dm/SsRS3KMA6oz6Kk/
A3Lz1s9uxmkLb5JqX9Gwvn1GUH3eiVhQgtv6ORCbedkKPp3iMtFJ+m5bImAEN5XXYo5t9cb5E5Wf
ZklQS0+1gnvxS/piphUZdGjkfFLUSbKPq7MULXEA2Gb2bs8lIfVjy//U+S5b977PvshP/GOutTCf
lSC95uLh0utmHUryjW6TOPqHPgQmo5mHJuQueTXReuzFsEThdoYyDFW+4TYKN+TLPt/eKNlySIkG
4ivtEwCoDTe0n4GgzzC3gisP3u8GM0k8rAlhzkD4PiR+q/r3g0E08o5BFo+MOVZhL5/cVQHIEfNt
zpo6EEqHyLHv6V+C+PveAoRZB9eZC/Ke1jGlcazMCBDqttmYDjWqDycTigcNkygCvcmKHAHIxQKH
V0WVf4kj9IIB/50xnnmHVcHt4m8o4SrNdlBQ1yGOD3ZSDrHj1BoK9U0dCH6sBT8c+JTzghq/vMgg
OrIr99QvRIBB2i6xs2UzvjviPfxRBClwWo6rTtzRtqexF68Zi16wS3TKs5ME3je4ypNyYpR5Fyxh
U8sW45CPuiB0cHCQiJa50En1h45wQi6U2SG+kFTAG6cyPSc8EWc5Gb/jrc3uDOhyy7fg5hGeOjje
5sq0R6PVvsBOkp23tnEJBkPDFSFTbbpklBPx0j4Q1oAHBhXYFTViAXndGtt9cgch7SFErHEXEXNA
POmAws/dsh6QOTBAcrvc880YhEod1wsamjnelcgj/cZnixu3XPqBmB+PB/cS+GK0Im1qtv2PdczJ
V7S+G7GcnFiXh5ZoNspLts9ZNgc1Orqj05IPH/rPjLtGgy99cRYOak9TfRVDqqBgezjRFpOPTswR
uxkCYcwaCJrNgJn0fbHoMfmlNMlFoxYHd1ZbMUOhcMpCHEBm3PBtzoKrR0l6tw/FsQho2BsLJryV
WawN1S0SRiQiHTabi6RAsXCfgjIXIzt3oqDCISc2q4tUcjPK9AvD3Ql0w3CiwzEoP/b0zKTsUp8S
RChEGSGCBmPiSmmTw/ojQRK4E7McMbgxzjMTo8LBhS/BNB3y7YFhuHa2g+X5cYvM7t5tSW0SxuOg
HI9Q7HH6WhkQKn1LjijKLk6K/n/qdobbWgGLOCk08G/j+nF4qsH0phqrHangLtiBM9k9gsiMDqg1
siENbklaWz5AaWBn8PsYQVmz6ZQg/FnZ83mewQKY8hVW+pc8OSRvHsEl81KuJs1Qii7pJz3B38dG
Q8WLWL7cI5l38YhsN0Zt/F6Op4k6Xnq+JqlO8QwuggWEHlszOw2sdwsxAj2kHsA36AiH32EVxTvX
f0fffOLXmMWEJ6hTN6pwSN2f3MvGjEKLvnPUUcG1cqnT6cV26qyUqIiQ4DLLzoixZ+KxKFyp06wH
XRiS42CJU02kwPgTMlDn4XbLrrcZ+iIgh6XXweata+/j3TLAJ2/aRf/CC5UIr628xqggUFSWJDUn
W5QZvJtncSYKStc0ITEKtUvB6+6A7xGjYlpi2p0bkIrokvuWTqmihF5soADpeYqxRsOkWkBNM5oi
PgUB1YZwkAKrOBXchbMUotDnENrMFDEkprIVhShxcUuHetb8R4B6x2J2nKVSoqJDs/a2CaJcRSEn
gD7aN7DfrgnWrC1g1oY1trjltY1gV04frYNC89RZDnZHopYCAFI61QIrD+hmmR+Vgg9ZuOBN9GL4
0xpX3ysqZleOcktAuyyngA44AqBoI/YUkZTJYeeOylbFsnen8WF/5ZoTYbWhZ4q0BIYO6mB4jHeL
aWBWCFhm9UfmXI+G4zE+IolovwxXsogWsYZYZU5zL9sudV7hxr9BDVV8w4r5T6WNB2wZnGNz8pxn
A2CMIhcaWyRhAqwJREIqMxA0cfVkuQsgild4+MWLyDuc6djWWnge0jitdXlYkmngsejQq2IACyTi
u9XD+CWk0m5xylmQvbp09Ta3JgLtcreu82EpfEgClVTf9erNMMkk3CZv7jwVaFJES6+W9b8MRSlA
pUIKukRxNEPMNTTOPqqA6g2xOoB0BU/Oogrx7QtL/o340BnvZe7IKYp0nuzFRDRkHirm+98ZQ6iW
NG9UJD+eI5ohELytV7v8OMFtRlzgfucgfM22MlZXBKTaC3+orU91Zg1xb9i4/58kym0x7NX6pkn6
hOAXzGQBs8eXdOb8PxFtn4bIgSVdsUwUMI7JMy3ug8eriegh5Z1Pycsydk0BUf/ig/CP0AJb/14K
h0gFYVzza5HZb7YHlcluF40DJUPoOO6oEUKWS+mydRM8DmlKfHKcQ5oFLIsY8ofhxlt0HLmUndIR
KEZf3kVs/WzjamJYqY/97fzuE/BJOVaiwihdW9ih1kCH4gTT3sW2tSmcLIfdX7lNAPKtbIDmKxce
dauBhsZTd8Qy2QJ72HEz3Nh7PRp5gc5CX1ZR/tF87UbcZF6taGoZVp9xfytN4RyftRZLJefzxti6
x0Vnl7UZVKXeeng7cYD1C2Pg9rfieYUvkgK6f75uyBUWD/bsLkIdBv5N6D/Cfh2rCm5z6w6a7fOU
23anZ3ITgxDn9VRvwQgzLFLn0xkCrf51mtbQKPFrPlx3YOmIZ/QIiLU3lD8fFscN3sWVVFXLkh5+
phmmHRdEiTfwNDE0mlOLTzZOs3hNwPDaoprsOgwj/Ax1LbSzRyKu/WuCwULABgP8Mj9S2iSvc6OY
n9IPEVDuylNUfxOzQNeMRTm6hAYGG9A8wHLT2mBxMKWOUAEz58EA9wkT6ijEZbvSPfA+zVDHUJq6
dioELVULrvPTHIKksX4bcd2KDIETLmExgf39BXfwoT+vak6dcacqnHpMkgLIOp3k+GG/Wn63kcpR
slGA0d7/zVnei0E9KDwKvG4ruC8sqPxGKUbwVQuc3IIsXBUzoJnggCodXgOG2a5qM4sNjXLnuWYM
aNirwbf2574ARl7rvnru7hVc+eUpTfpvwzA2ax34mwXj4t4YmrpR6vp6VvJNoXRekSwLY/NrhVBq
/xWOs7W5N5u/iSElzvz/97UtmgVQS/yHdNTGqe+K8Fnoqgf+gIRLLNR+zNAoot568tU+nfz8zMrV
amxVO+A9HGTSIFmR0v9tjdh4k2IPTxf8n2jXBhE1AFmpjzgzLXZSXI61UR+ZMJ6gKB9IrQuDbuJe
7A4qpoJAYF5ideO/AICAQnbf9ZBHmq4GC83YrnsA7f/x/cHJhDd8/TUER0RL2VDnN67DU2Pp1C0O
jHT6cARMH2X0EkYkLi11b3e1rghF4nT6VN+KUNS4ejptLnRxcjtZZA3D/JETn9kYy5XTAfBuwlYj
pmmvk52V+wX6vXYuYMsWiRH/ngRzawHvUs+DRaQ/maVL6+5I7Q+lSW86+K0sFngfIHFlEfn3hW8O
YT2uJS52h5YMbfebs/y5rPyzgENOpNUsgJj7ApsZkb2j7MvD+az3Yp6X0NL46gy2CDvdMB0ha3qE
gPzO4fvQeMivHScTzCHvagpAIZycrscQ9bzAz5oWzPkv18NIsh7uOY0tDCfwaKh7t/0gigmpHYNm
FgUiGwBNdAItwlWNOwbaQRqvlumDsjuMmas9oEHbgqaqF/Wz2j/jTnHsA3xMOyGlvxS7BP3O5CZI
S/XQ1M4+KHQc5Hps4TG2V1PkMP/heMx1bVehexFOcixJOWVhFBQF9djc7dYvmbjxacRmeacMMPTB
4Poms/jp53DOw9ygkMFy89sI+Hqe5/uj2NMmfJXCuKRe6w5j1B4CfS9Egh/OJEchYPpVm3D47fys
0lmFuc7iVKc0z8QyqdOl9P23XA0PhLNYgYR2F3Z2xzKKqiygZWYdQSB7mYe64jmpauKAHJw1OKxB
lOcsiZuiVoX5zgOXjSh4781UmxVjfOCMxO+ePR1QBBdaIk0MfLlA3ZJBsWFf9Ape8wqfg65fhnT4
K1w5lflmznAqXl8KcButbsG/rOFf4SglRGVwDcjmh20JW/ODx//YCe1X2LoeZobAT+hhVBW0E5qv
7HFL2g+UubpCAkwgFp7I3zThxWAfdiyyKxKVgD451M3wDLqhaeFjCOr76ypJcSKTUgVzcbz0PkfJ
Rx4loliDYiKbPdlLUuRl/uddEOo1ilcdyc9PsX+umWfu9EiThUQGOy/ssoN08CMIRcpRjCdBs1jT
AOWWG68ZhtHuW80yJW1PUl1ARaikLpixNXnVQjZjGFpzH4+HUQjttBKzxkdKQBc+ZVYDiODlw7lo
tvsdgZpkHeISPW7QO2qvJWWxNMNI5tV57fu+V3ZgY65H95giYfm0BowshSVMd73Fq8FqDsqjFCq1
wVASqth+BidlCgqOC2H91iMxfu2e6EMiAmT1HpYFttk0i/TsT9ZPZa78o4S6lEtNHXg+1jReiifi
Uc4YVvwmL7C50dJe6RXvmtryBBe8F81Gy5KDSCwXOP1QLo0ai6srua5tHDp+zu0WIwxYhSrEA9sT
ZmSC5LbvCzOuel/GybUz7aQp4CvrSDe6GVhE+pGar8CBOS+CxsUF/ElRCBz3juHlGxQQ
`protect end_protected
